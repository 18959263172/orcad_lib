-- "$Header: act3.vhd@@/main/4 $"
-- Actel Vital 95 library for R299 release.
library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;

package COMPONENTS is

constant DefaultTimingChecksOn : Boolean := True;
constant DefaultXGenerationOn : Boolean := False;
constant DefaultXon : Boolean := False;
constant DefaultMsgOn : Boolean := True;

component AND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND5B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO10
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO11
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO5A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO6
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO6A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO7
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO8
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO9
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BBHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BBHSA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_IDE_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BBLSA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_IDE_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BBUFTH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BBUFTL
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BIBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BIECTH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BIECTL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns); 	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BIEPTH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns); 	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BIEPTL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns); 	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BRECTH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BRECTL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BREPTH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BREPTL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component BUFA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BUFF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CLKBIBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CLKBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CLKINT
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CM7
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CM8
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S01_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S00_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CS1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CS2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CY2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CY2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component DECETH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component DECETL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component DEPETH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component DEPETL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component DF1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DF1A_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DF1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DF1C_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFC1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1A_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1D_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFC1G
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFE
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1C_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFEA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFEA_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM1C_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM3E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM6A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM6B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM7A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM7B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM8A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S00_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S00_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S01_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S01_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S00                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S01                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM8B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S00_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S00_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S01_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S01_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFMA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFMA_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFMB
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFME1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1A_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFP1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1D_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFP1F
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFP1G
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFPC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFPC_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFPCA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFPCA_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DL1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DL2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DL2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL2D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLC1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLC1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLC1F
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLC1G
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLCA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLE2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLEA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLEB
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLEC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM8A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S00_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S01_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S00_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S00_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S01_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S01_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S00                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S01                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM8B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S00_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S01_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S00_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S00_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S01_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S01_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S00                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S01                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLMA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLME1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_A_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_A_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_B_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_B_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_S_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLP1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component FA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
end component; 

component FA1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
end component; 

component FA2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
end component; 

component FECTH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
                tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);        -- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component FECTL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
                tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);        -- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component FECTMH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component FECTML
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component FEPTH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component FEPTL
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component FEPTMH
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component FEPTML
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	--
end component; 

component GAND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GMX4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GNAND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GND
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '0');
end component; 

component GNOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GXOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component HA1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component HA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component HA1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component HA1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component HCLKBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component IBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component INBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component INV
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component INVA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component IOCLKBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component IODFE
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component IODFEC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component IODFEP
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component IOPCLBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component IREC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_IDE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_IDE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      PAD                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component IREP
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_IDE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_IDE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      PAD                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component MAJ3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MXC1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MXT
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0B_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0A_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0A                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0B                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0A                            :	in    STD_ULOGIC;
      S0B                            :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND5C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR5C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA5
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OBHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OBUFTH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OBUFTL
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR5B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component ORECTH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component ORECTL
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OREPTH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OREPTL
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OUTBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component TBHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component TF1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component TF1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component TRIBUFF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component VCC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '1');
end component; 

component XA1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XNOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XO1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XO1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

end COMPONENTS;

----------------------------------------------------------------
-- 
-- 
----------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;
use IEEE.VITAL_Primitives.all;

package VTABLES is

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DF1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   CONSTANT DF1A_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  H ),
    ( L,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ));

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ));

   CONSTANT DFC1E_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  H,  x,  L ),
    ( L,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( x,  L,  x,  x,  x,  H ),
    ( x,  H,  x,  L,  x,  S ));

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFE3A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  H,  H,  x,  L ));

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ));

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ));

   CONSTANT DFM4C_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  H,  H,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  H,  x,  L ));

   CONSTANT DFM6A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  x,  L ));

   CONSTANT DFM7A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  L,  H,  x,  L ));

   CONSTANT DFM8A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  H,  H,  x,  L ));

   CONSTANT DFME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H,  L,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  H,  x,  H,  L,  H,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ));

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ));

   CONSTANT DFP1C_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  L,  x,  H ),
    ( L,  H,  H,  x,  x,  L ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ));

   CONSTANT DFP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  H,  H,  x,  L ));

   CONSTANT DFPC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ));

   CONSTANT DL1_Q_tab : VitalStateTableType := (
    ( L,  H,  x,  L ),
    ( H,  H,  x,  H ),
    ( x,  L,  x,  S ));

   CONSTANT DL1A_QN_tab : VitalStateTableType := (
    ( L,  H,  x,  H ),
    ( H,  H,  x,  L ),
    ( x,  L,  x,  S ));

   CONSTANT DL1B_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  L ),
    ( L,  H,  x,  H ),
    ( H,  x,  x,  S ));

   CONSTANT DL1C_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  H ),
    ( L,  H,  x,  L ),
    ( H,  x,  x,  S ));

   CONSTANT DL2A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  L,  x,  S ),
    ( H,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  H,  x,  L ));

   CONSTANT DL2B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  H,  x,  x,  S ),
    ( L,  x,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  L,  x,  H ));

   CONSTANT DL2C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  x,  H ),
    ( H,  H,  x,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  H ),
    ( x,  L,  L,  L,  x,  L ));

   CONSTANT DL2D_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  x,  L,  x,  S ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  H,  x,  H ));

   CONSTANT DLC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  L,  H,  x,  L ));

   CONSTANT DLC1_Q_tab : VitalStateTableType := (
    ( L,  H,  x,  x,  L ),
    ( H,  H,  L,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  L ));

   CONSTANT DLC1A_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  L ),
    ( L,  H,  L,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  L ));

   CONSTANT DLC1F_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( L,  x,  L,  x,  S ),
    ( H,  x,  x,  x,  H ),
    ( x,  L,  H,  x,  H ));

   CONSTANT DLC1G_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H ),
    ( H,  L,  x,  x,  S ),
    ( x,  H,  x,  x,  H ));

   CONSTANT DLCA_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  L,  x,  L ));

   CONSTANT DLE_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( x,  L,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   CONSTANT DLE1D_QN_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H ),
    ( L,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   CONSTANT DLE2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  L ));

   CONSTANT DLE2C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ));

   CONSTANT DLE3B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  H ));

   CONSTANT DLE3C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  H,  x,  S ),
    ( x,  H,  x,  H,  x,  S ),
    ( x,  x,  x,  L,  x,  H ));

   CONSTANT DLEC_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   CONSTANT DLM_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  H,  x,  H ),
    ( x,  L,  L,  H,  x,  L ),
    ( x,  H,  L,  H,  x,  H ),
    ( x,  x,  x,  L,  x,  S ));

   CONSTANT DLM2_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  x,  L ),
    ( x,  x,  L,  L,  H,  x,  L ));

   CONSTANT DLM2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  x,  L ));

   CONSTANT DLM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DLM3A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ));

   CONSTANT DLM4_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DLM4A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  S ));

   CONSTANT DLM8A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  H,  H,  H,  H,  x,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  H,  x,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  H,  x,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  x,  x,  x,  L,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  x,  x,  x,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  L,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  x,  H,  x,  H,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  H,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  x,  H,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  H,  H,  L,  L,  x,  x,  H,  x,  H ),
    ( H,  x,  x,  H,  x,  L,  L,  L,  x,  H,  x,  H ),
    ( H,  x,  x,  H,  x,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  L,  L,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  H,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  x,  H,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  x,  L,  x,  x,  H,  x,  H,  H,  H,  x,  L ),
    ( x,  x,  L,  x,  x,  x,  H,  H,  H,  H,  x,  L ),
    ( x,  x,  x,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  x,  x,  x,  L,  L,  L,  H,  H,  H,  x,  L ));

   CONSTANT DLM8B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  x,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  x,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  L,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  x,  L,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  L,  x,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  x,  L,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  L,  x,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  x,  L,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  x,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  L,  x,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  x,  L,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  x,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  x,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  x,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  x,  L,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  x,  L,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  x,  L,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  x,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  L,  x,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  x,  L,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  H,  x,  L ));

   CONSTANT DLMA_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  x,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L ),
    ( L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  S ));

   CONSTANT DLME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  H,  H,  x,  x,  H ),
    ( L,  L,  H,  x,  H,  x,  H ),
    ( L,  L,  x,  L,  L,  x,  L ),
    ( L,  L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  x,  x,  S ));

   CONSTANT DLP1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  H,  x,  x,  H ));

   CONSTANT DLP1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  H ));

   CONSTANT DLP1B_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  x,  x,  H ),
    ( x,  H,  L,  x,  S ));

   CONSTANT DLP1C_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  H,  x,  S ),
    ( x,  x,  L,  x,  H ));

   CONSTANT DLP1D_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  H,  H,  x,  L ));

   CONSTANT DLP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  H,  x,  L ));

   CONSTANT IODFEP_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  x,  H ),
    ( x,  x,  x,  x,  H,  L,  x,  S ));

   CONSTANT TF1A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( x,  L,  H,  H,  H,  x,  L ));


end VTABLES;

---- end of VITAL tables library ----
----- CELL AND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND2 : entity is TRUE;
end AND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND2_VITAL of AND2 is
   for VITAL_ACT
   end for;
end CFG_AND2_VITAL;


----- CELL AND2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND2A : entity is TRUE;
end AND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND2A_VITAL of AND2A is
   for VITAL_ACT
   end for;
end CFG_AND2A_VITAL;


----- CELL AND2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND2B : entity is TRUE;
end AND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND2B_VITAL of AND2B is
   for VITAL_ACT
   end for;
end CFG_AND2B_VITAL;


----- CELL AND3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3 : entity is TRUE;
end AND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND (A_ipd) AND (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3_VITAL of AND3 is
   for VITAL_ACT
   end for;
end CFG_AND3_VITAL;


----- CELL AND3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3A : entity is TRUE;
end AND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND ((NOT A_ipd)) AND (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3A_VITAL of AND3A is
   for VITAL_ACT
   end for;
end CFG_AND3A_VITAL;


----- CELL AND3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3B : entity is TRUE;
end AND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3B_VITAL of AND3B is
   for VITAL_ACT
   end for;
end CFG_AND3B_VITAL;


----- CELL AND3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3C : entity is TRUE;
end AND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3C_VITAL of AND3C is
   for VITAL_ACT
   end for;
end CFG_AND3C_VITAL;


----- CELL AND4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4 : entity is TRUE;
end AND4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND (A_ipd) AND (C_ipd) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4_VITAL of AND4 is
   for VITAL_ACT
   end for;
end CFG_AND4_VITAL;


----- CELL AND4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4A : entity is TRUE;
end AND4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4A_VITAL of AND4A is
   for VITAL_ACT
   end for;
end CFG_AND4A_VITAL;


----- CELL AND4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4B : entity is TRUE;
end AND4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4B_VITAL of AND4B is
   for VITAL_ACT
   end for;
end CFG_AND4B_VITAL;


----- CELL AND4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4C : entity is TRUE;
end AND4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4C_VITAL of AND4C is
   for VITAL_ACT
   end for;
end CFG_AND4C_VITAL;


----- CELL AND4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4D : entity is TRUE;
end AND4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND ((NOT D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4D_VITAL of AND4D is
   for VITAL_ACT
   end for;
end CFG_AND4D_VITAL;


----- CELL AND5B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND5B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND5B : entity is TRUE;
end AND5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AND5B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd) AND (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND5B_VITAL of AND5B is
   for VITAL_ACT
   end for;
end CFG_AND5B_VITAL;


----- CELL AO1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1 : entity is TRUE;
end AO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1_VITAL of AO1 is
   for VITAL_ACT
   end for;
end CFG_AO1_VITAL;


----- CELL AO10 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO10 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO10 : entity is TRUE;
end AO10;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO10 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((E_ipd) OR (D_ipd)) AND ((C_ipd) OR ((B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO10_VITAL of AO10 is
   for VITAL_ACT
   end for;
end CFG_AO10_VITAL;


----- CELL AO11 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO11 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO11 : entity is TRUE;
end AO11;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO11 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((C_ipd) AND ((B_ipd) OR (A_ipd))) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO11_VITAL of AO11 is
   for VITAL_ACT
   end for;
end CFG_AO11_VITAL;


----- CELL AO1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1A : entity is TRUE;
end AO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1A_VITAL of AO1A is
   for VITAL_ACT
   end for;
end CFG_AO1A_VITAL;


----- CELL AO1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1B : entity is TRUE;
end AO1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1B_VITAL of AO1B is
   for VITAL_ACT
   end for;
end CFG_AO1B_VITAL;


----- CELL AO1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1C : entity is TRUE;
end AO1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1C_VITAL of AO1C is
   for VITAL_ACT
   end for;
end CFG_AO1C_VITAL;


----- CELL AO1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1D : entity is TRUE;
end AO1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1D_VITAL of AO1D is
   for VITAL_ACT
   end for;
end CFG_AO1D_VITAL;


----- CELL AO1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1E : entity is TRUE;
end AO1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1E_VITAL of AO1E is
   for VITAL_ACT
   end for;
end CFG_AO1E_VITAL;


----- CELL AO2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2 : entity is TRUE;
end AO2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND (A_ipd)) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2_VITAL of AO2 is
   for VITAL_ACT
   end for;
end CFG_AO2_VITAL;


----- CELL AO2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2A : entity is TRUE;
end AO2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2A_VITAL of AO2A is
   for VITAL_ACT
   end for;
end CFG_AO2A_VITAL;


----- CELL AO2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2B : entity is TRUE;
end AO2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2B_VITAL of AO2B is
   for VITAL_ACT
   end for;
end CFG_AO2B_VITAL;


----- CELL AO2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2C : entity is TRUE;
end AO2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2C_VITAL of AO2C is
   for VITAL_ACT
   end for;
end CFG_AO2C_VITAL;


----- CELL AO2D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2D : entity is TRUE;
end AO2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO2D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2D_VITAL of AO2D is
   for VITAL_ACT
   end for;
end CFG_AO2D_VITAL;


----- CELL AO2E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2E : entity is TRUE;
end AO2E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO2E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd))) OR ((NOT D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2E_VITAL of AO2E is
   for VITAL_ACT
   end for;
end CFG_AO2E_VITAL;


----- CELL AO3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3 : entity is TRUE;
end AO3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR ((B_ipd) AND ((NOT A_ipd)) AND (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3_VITAL of AO3 is
   for VITAL_ACT
   end for;
end CFG_AO3_VITAL;


----- CELL AO3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3A : entity is TRUE;
end AO3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR ((B_ipd) AND (A_ipd) AND (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3A_VITAL of AO3A is
   for VITAL_ACT
   end for;
end CFG_AO3A_VITAL;


----- CELL AO3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3B : entity is TRUE;
end AO3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3B_VITAL of AO3B is
   for VITAL_ACT
   end for;
end CFG_AO3B_VITAL;


----- CELL AO3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3C : entity is TRUE;
end AO3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (D_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3C_VITAL of AO3C is
   for VITAL_ACT
   end for;
end CFG_AO3C_VITAL;


----- CELL AO4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO4A : entity is TRUE;
end AO4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of AO4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((C_ipd) AND (A_ipd) AND (D_ipd)) OR ((B_ipd) AND ((NOT A_ipd)) AND
         (C_ipd)) OR ((C_ipd) AND (B_ipd) AND (D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO4A_VITAL of AO4A is
   for VITAL_ACT
   end for;
end CFG_AO4A_VITAL;


----- CELL AO5A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO5A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO5A : entity is TRUE;
end AO5A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of AO5A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((C_ipd) AND (A_ipd)) OR ((B_ipd) AND ((NOT A_ipd))) OR ((C_ipd) AND (B_ipd)) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO5A_VITAL of AO5A is
   for VITAL_ACT
   end for;
end CFG_AO5A_VITAL;


----- CELL AO6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO6 : entity is TRUE;
end AO6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO6 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) AND (C_ipd)) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO6_VITAL of AO6 is
   for VITAL_ACT
   end for;
end CFG_AO6_VITAL;


----- CELL AO6A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO6A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO6A : entity is TRUE;
end AO6A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO6A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (((NOT D_ipd)) AND (C_ipd)) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO6A_VITAL of AO6A is
   for VITAL_ACT
   end for;
end CFG_AO6A_VITAL;


----- CELL AO7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO7 : entity is TRUE;
end AO7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO7 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR ((B_ipd) AND (A_ipd) AND (C_ipd)) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO7_VITAL of AO7 is
   for VITAL_ACT
   end for;
end CFG_AO7_VITAL;


----- CELL AO8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO8 : entity is TRUE;
end AO8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO8 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (((NOT D_ipd)) AND ((NOT C_ipd))) OR ((B_ipd) AND (A_ipd)) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO8_VITAL of AO8 is
   for VITAL_ACT
   end for;
end CFG_AO8_VITAL;


----- CELL AO9 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO9 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO9 : entity is TRUE;
end AO9;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AO9 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND (A_ipd)) OR (D_ipd) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO9_VITAL of AO9 is
   for VITAL_ACT
   end for;
end CFG_AO9_VITAL;


----- CELL AOI1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1 : entity is TRUE;
end AOI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1_VITAL of AOI1 is
   for VITAL_ACT
   end for;
end CFG_AOI1_VITAL;


----- CELL AOI1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1A : entity is TRUE;
end AOI1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR ((B_ipd) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1A_VITAL of AOI1A is
   for VITAL_ACT
   end for;
end CFG_AOI1A_VITAL;


----- CELL AOI1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1B : entity is TRUE;
end AOI1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT C_ipd)) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1B_VITAL of AOI1B is
   for VITAL_ACT
   end for;
end CFG_AOI1B_VITAL;


----- CELL AOI1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1C : entity is TRUE;
end AOI1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1C_VITAL of AOI1C is
   for VITAL_ACT
   end for;
end CFG_AOI1C_VITAL;


----- CELL AOI1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1D : entity is TRUE;
end AOI1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1D_VITAL of AOI1D is
   for VITAL_ACT
   end for;
end CFG_AOI1D_VITAL;


----- CELL AOI2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI2A : entity is TRUE;
end AOI2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI2A_VITAL of AOI2A is
   for VITAL_ACT
   end for;
end CFG_AOI2A_VITAL;


----- CELL AOI2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI2B : entity is TRUE;
end AOI2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT C_ipd)) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI2B_VITAL of AOI2B is
   for VITAL_ACT
   end for;
end CFG_AOI2B_VITAL;


----- CELL AOI3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI3A : entity is TRUE;
end AOI3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (A_ipd)) AND ((B_ipd) OR (A_ipd) OR (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI3A_VITAL of AOI3A is
   for VITAL_ACT
   end for;
end CFG_AOI3A_VITAL;


----- CELL AOI4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI4 : entity is TRUE;
end AOI4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((D_ipd) AND (C_ipd)) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI4_VITAL of AOI4 is
   for VITAL_ACT
   end for;
end CFG_AOI4_VITAL;


----- CELL AOI4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI4A : entity is TRUE;
end AOI4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AOI4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((D_ipd) AND ((NOT C_ipd))) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI4A_VITAL of AOI4A is
   for VITAL_ACT
   end for;
end CFG_AOI4A_VITAL;


----- CELL AX1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1 : entity is TRUE;
end AX1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AX1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) XOR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1_VITAL of AX1 is
   for VITAL_ACT
   end for;
end CFG_AX1_VITAL;


----- CELL AX1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1A : entity is TRUE;
end AX1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AX1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) XOR ((B_ipd) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1A_VITAL of AX1A is
   for VITAL_ACT
   end for;
end CFG_AX1A_VITAL;


----- CELL AX1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1B : entity is TRUE;
end AX1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AX1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) XOR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1B_VITAL of AX1B is
   for VITAL_ACT
   end for;
end CFG_AX1B_VITAL;


----- CELL AX1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1C : entity is TRUE;
end AX1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of AX1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) XOR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1C_VITAL of AX1C is
   for VITAL_ACT
   end for;
end CFG_AX1C_VITAL;


----- CELL BBHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BBHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BBHS : entity is TRUE;
end BBHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BBHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BBHS_VITAL of BBHS is
   for VITAL_ACT
   end for;
end CFG_BBHS_VITAL;


----- CELL BBHSA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BBHSA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_IDE_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BBHSA : entity is TRUE;
end BBHSA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BBHSA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IDE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (IDE_ipd, IDE, tipd_IDE);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, IDE_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := (PAD_ipd) AND (IDE_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (IDE_ipd'last_event, tpd_IDE_Y, TRUE),
                 1 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BBHSA_VITAL of BBHSA is
   for VITAL_ACT
   end for;
end CFG_BBHSA_VITAL;


----- CELL BBLSA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BBLSA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_IDE_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BBLSA : entity is TRUE;
end BBLSA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BBLSA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IDE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (IDE_ipd, IDE, tipd_IDE);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, IDE_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := (PAD_ipd) AND (IDE_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (IDE_ipd'last_event, tpd_IDE_Y, TRUE),
                 1 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BBLSA_VITAL of BBLSA is
   for VITAL_ACT
   end for;
end CFG_BBLSA_VITAL;


----- CELL BBUFTH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BBUFTH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BBUFTH : entity is TRUE;
end BBUFTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BBUFTH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BBUFTH_VITAL of BBUFTH is
   for VITAL_ACT
   end for;
end CFG_BBUFTH_VITAL;


----- CELL BBUFTL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BBUFTL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BBUFTL : entity is TRUE;
end BBUFTL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BBUFTL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BBUFTL_VITAL of BBUFTL is
   for VITAL_ACT
   end for;
end CFG_BBUFTL_VITAL;


----- CELL BIBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BIBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BIBUF : entity is TRUE;
end BIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BIBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BIBUF_VITAL of BIBUF is
   for VITAL_ACT
   end for;
end CFG_BIBUF_VITAL;


















----- CELL BIECTH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BIECTH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BIECTH : ENTITY IS TRUE;
	--
end BIECTH;

ARCHITECTURE VITAL_ACT OF BIECTH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  BIECTH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  BIECTH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BIECTH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_BIECTH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : BIECTH_TAB Declaration
		CONSTANT  BIECTH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
                --Vio, Clr, Clk,   d,   e, prev, next 
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : BIECTH_TAB
		VitalStateTable (
				StateTable         => BIECTH_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => BIECTH_TAB_Result,
				PreviousDataIn     => PrevData_BIECTH_TAB
		);	--End VitalStateTable
		BIECTH_TABStateReg(0)     := BIECTH_TAB_Result(2);
		Q_zd                      := BIECTH_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => D_ipd, enable => (NOT E_ipd));
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;


		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => D_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_D_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BIECTH_VITAL of BIECTH is
   for VITAL_ACT
   end for;
end CFG_BIECTH_VITAL;
----- CELL BIECTL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BIECTL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns); 	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BIECTL : ENTITY IS TRUE;
	--
end BIECTL;

ARCHITECTURE VITAL_ACT OF BIECTL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  BIECTL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  BIECTL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BIECTL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_BIECTL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : BIECTL_TAB Declaration
		CONSTANT  BIECTL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
                --Vio, Clr, Clk,   d,   e, prev, next 
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : BIECTL_TAB
		VitalStateTable (
				StateTable         => BIECTL_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => BIECTL_TAB_Result,
				PreviousDataIn     => PrevData_BIECTL_TAB
		);	--End VitalStateTable
		BIECTL_TABStateReg(0)     := BIECTL_TAB_Result(2);
		Q_zd                      := BIECTL_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => D_ipd, enable => (NOT E_ipd));
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;


		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => D_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_D_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BIECTL_VITAL of BIECTL is
   for VITAL_ACT
   end for;
end CFG_BIECTL_VITAL;
----- CELL BIEPTH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BIEPTH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns); 	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BIEPTH : ENTITY IS TRUE;
	--
end BIEPTH;

ARCHITECTURE VITAL_ACT OF BIEPTH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  BIEPTH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  BIEPTH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BIEPTH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 5);
		--VARIABLE  PrevData_BIEPTH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_BIEPTH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : BIEPTH_TAB Declaration
		CONSTANT  BIEPTH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
--          Violation, IOPCL, CLK, D, ODE
		( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : BIEPTH_TAB
		VitalStateTable (
				StateTable         => BIEPTH_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => BIEPTH_TAB_Result,
				PreviousDataIn     => PrevData_BIEPTH_TAB
		);	--End VitalStateTable
		BIEPTH_TABStateReg(0)     := BIEPTH_TAB_Result(2);
		Q_zd                      := BIEPTH_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => D_ipd, enable => (NOT E_ipd));
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => D_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_D_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BIEPTH_VITAL of BIEPTH is
   for VITAL_ACT
   end for;
end CFG_BIEPTH_VITAL;
----- CELL BIEPTL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BIEPTL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_D_PAD            : VitalDelayType01 := (1.000 ns, 1.000 ns); 	-- Path delay from input D to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BIEPTL : ENTITY IS TRUE;
	--
end BIEPTL;

ARCHITECTURE VITAL_ACT OF BIEPTL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  BIEPTL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  BIEPTL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BIEPTL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 5);
		--VARIABLE  PrevData_BIEPTL_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_BIEPTL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : BIEPTL_TAB Declaration
		CONSTANT  BIEPTL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
--          Violation, IOPCL, CLK, D, ODE
		( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : BIEPTL_TAB
		VitalStateTable (
				StateTable         => BIEPTL_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => BIEPTL_TAB_Result,
				PreviousDataIn     => PrevData_BIEPTL_TAB
		);	--End VitalStateTable
		BIEPTL_TABStateReg(0)     := BIEPTL_TAB_Result(2);
		Q_zd                      := BIEPTL_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => D_ipd, enable => (NOT E_ipd));
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => D_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_D_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BIEPTL_VITAL of BIEPTL is
   for VITAL_ACT
   end for;
end CFG_BIEPTL_VITAL;
----- CELL BRECTH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BRECTH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BRECTH : ENTITY IS TRUE;
	--
end BRECTH;

ARCHITECTURE VITAL_ACT OF BRECTH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  BRECTH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  BRECTH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BRECTH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_BRECTH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_BRECTH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : BRECTH_TAB Declaration
		CONSTANT  BRECTH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : BRECTH_TAB
		VitalStateTable (
				StateTable         => BRECTH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => BRECTH_TAB_Result,
				PreviousDataIn     => PrevData_BRECTH_TAB
		);	--End VitalStateTable
		BRECTH_TABStateReg(0)     := BRECTH_TAB_Result(2);
		IQ(0)                     := BRECTH_TAB_Result(1);
		Y_zd                      := TO_X01(PAD_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BRECTH_VITAL of BRECTH is
   for VITAL_ACT
   end for;
end CFG_BRECTH_VITAL;
----- CELL BRECTL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BRECTL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BRECTL : ENTITY IS TRUE;
	--
end BRECTL;

ARCHITECTURE VITAL_ACT OF BRECTL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  BRECTL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  BRECTL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BRECTL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_BRECTL_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_BRECTL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : BRECTL_TAB Declaration
		CONSTANT  BRECTL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : BRECTL_TAB
		VitalStateTable (
				StateTable         => BRECTL_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => BRECTL_TAB_Result,
				PreviousDataIn     => PrevData_BRECTL_TAB
		);	--End VitalStateTable
		BRECTL_TABStateReg(0)     := BRECTL_TAB_Result(2);
		IQ(0)                     := BRECTL_TAB_Result(1);
		Y_zd                      := TO_X01(PAD_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BRECTL_VITAL of BRECTL is
   for VITAL_ACT
   end for;
end CFG_BRECTL_VITAL;
----- CELL BREPTH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BREPTH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BREPTH : ENTITY IS TRUE;
	--
end BREPTH;

ARCHITECTURE VITAL_ACT OF BREPTH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  BREPTH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  BREPTH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BREPTH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_BREPTH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_BREPTH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : BREPTH_TAB Declaration
		CONSTANT  BREPTH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : BREPTH_TAB
		VitalStateTable (
				StateTable         => BREPTH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => BREPTH_TAB_Result,
				PreviousDataIn     => PrevData_BREPTH_TAB
		);	--End VitalStateTable
		BREPTH_TABStateReg(0)     := BREPTH_TAB_Result(2);
		IQ(0)                     := BREPTH_TAB_Result(1);
		Y_zd                      := TO_X01(PAD_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BREPTH_VITAL of BREPTH is
   for VITAL_ACT
   end for;
end CFG_BREPTH_VITAL;
----- CELL BREPTL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity BREPTL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF BREPTL : ENTITY IS TRUE;
	--
end BREPTL;

ARCHITECTURE VITAL_ACT OF BREPTL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  BREPTL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  BREPTL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  BREPTL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_BREPTL_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_BREPTL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : BREPTL_TAB Declaration
		CONSTANT  BREPTL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : BREPTL_TAB
		VitalStateTable (
				StateTable         => BREPTL_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => BREPTL_TAB_Result,
				PreviousDataIn     => PrevData_BREPTL_TAB
		);	--End VitalStateTable
		BREPTL_TABStateReg(0)     := BREPTL_TAB_Result(2);
		IQ(0)                     := BREPTL_TAB_Result(1);
		Y_zd                      := TO_X01(PAD_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_BREPTL_VITAL of BREPTL is
   for VITAL_ACT
   end for;
end CFG_BREPTL_VITAL;
----- CELL BUFA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFA : entity is TRUE;
end BUFA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BUFA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BUFA_VITAL of BUFA is
   for VITAL_ACT
   end for;
end CFG_BUFA_VITAL;


----- CELL BUFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFF : entity is TRUE;
end BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of BUFF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BUFF_VITAL of BUFF is
   for VITAL_ACT
   end for;
end CFG_BUFF_VITAL;


----- CELL CLKBIBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBIBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBIBUF : entity is TRUE;
end CLKBIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of CLKBIBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBIBUF_VITAL of CLKBIBUF is
   for VITAL_ACT
   end for;
end CFG_CLKBIBUF_VITAL;


----- CELL CLKBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBUF : entity is TRUE;
end CLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of CLKBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBUF_VITAL of CLKBUF is
   for VITAL_ACT
   end for;
end CFG_CLKBUF_VITAL;


----- CELL CLKINT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKINT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKINT : entity is TRUE;
end CLKINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of CLKINT is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKINT_VITAL of CLKINT is
   for VITAL_ACT
   end for;
end CFG_CLKINT_VITAL;


----- CELL CM7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CM7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CM7 : entity is TRUE;
end CM7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CM7 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE OR_Out, MUX1_Out, MUX2_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- (((S11_ipd) OR (S10_ipd)) AND (((S0_ipd) AND (D3_ipd)) OR (((NOT
      --   S0_ipd)) AND (D2_ipd)))) OR (((NOT ((S11_ipd) OR (S10_ipd)))) AND
      --   (((S0_ipd) AND (D1_ipd)) OR (((NOT S0_ipd)) AND (D0_ipd))));
      OR_Out := VitalOR2(S10_ipd, S11_ipd);
      MUX1_Out := VitalMUX2(D1_ipd, D0_ipd, S0_ipd);
      MUX2_Out := VitalMUX2(D3_ipd, D2_ipd, S0_ipd);
      Y_zd := VitalMUX2(MUX2_Out, MUX1_Out, OR_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S11_ipd'last_event, tpd_S11_Y, TRUE),
                 1 => (S10_ipd'last_event, tpd_S10_Y, TRUE),
                 2 => (S0_ipd'last_event, tpd_S0_Y, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 4 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 5 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 6 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CM7_VITAL of CM7 is
   for VITAL_ACT
   end for;
end CFG_CM7_VITAL;


----- CELL CM8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CM8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S01_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S00_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CM8 : entity is TRUE;
end CM8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CM8 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S00_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S01_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S00_ipd, S00, tipd_S00);
   VitalWireDelay (S01_ipd, S01, tipd_S01);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S00_ipd, S01_ipd, S10_ipd, S11_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE AND_Out, OR_Out, MUX1_Out, MUX2_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- (((S11_ipd) OR (S10_ipd)) AND (((S01_ipd) AND (S00_ipd) AND (D3_ipd))
      --   OR (((NOT ((S01_ipd) AND (S00_ipd)))) AND (D2_ipd)))) OR (((NOT
      --   ((S11_ipd) OR (S10_ipd)))) AND (((S01_ipd) AND (S00_ipd) AND
      --   (D1_ipd)) OR (((NOT ((S01_ipd) AND (S00_ipd)))) AND (D0_ipd))));
      AND_Out := VitalAND2(S00_ipd, S01_ipd);
      OR_Out := VitalOR2(S10_ipd, S11_ipd);
      MUX1_Out := VitalMUX2(D1_ipd, D0_ipd, AND_Out);
      MUX2_Out := VitalMUX2(D3_ipd, D2_ipd, AND_Out);
      Y_zd := VitalMUX2(MUX2_Out, MUX1_Out, OR_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S11_ipd'last_event, tpd_S11_Y, TRUE),
                 1 => (S10_ipd'last_event, tpd_S10_Y, TRUE),
                 2 => (S01_ipd'last_event, tpd_S01_Y, TRUE),
                 3 => (S00_ipd'last_event, tpd_S00_Y, TRUE),
                 4 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 5 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 6 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 7 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CM8_VITAL of CM8 is
   for VITAL_ACT
   end for;
end CFG_CM8_VITAL;


----- CELL CS1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CS1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CS1 : entity is TRUE;
end CS1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CS1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE AND_Out, OR_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((((B_ipd) AND (S_ipd)) OR (A_ipd)) AND (D_ipd)) OR ((C_ipd) AND
      --   ((NOT (((B_ipd) AND (S_ipd)) OR (A_ipd)))));
      AND_Out := VitalAND2(B_ipd, S_ipd);
      OR_Out := VitalOR2(A_ipd, AND_Out);
      Y_zd := VitalMUX2(D_ipd, C_ipd, OR_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CS1_VITAL of CS1 is
   for VITAL_ACT
   end for;
end CFG_CS1_VITAL;


----- CELL CS2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CS2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CS2 : entity is TRUE;
end CS2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CS2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE AND_Out, OR_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((B_ipd) AND ((S_ipd) OR (A_ipd)) AND (D_ipd)) OR ((C_ipd) AND ((NOT
      --   ((B_ipd) AND ((S_ipd) OR (A_ipd))))));
      OR_Out := VitalOR2(A_ipd, S_ipd);
      AND_Out := VitalAND2(B_ipd, OR_Out);
      Y_zd := VitalMUX2(D_ipd, C_ipd, AND_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CS2_VITAL of CS2 is
   for VITAL_ACT
   end for;
end CFG_CS2_VITAL;


----- CELL CY2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CY2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CY2A : entity is TRUE;
end CY2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of CY2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B0_ipd, B0, tipd_B0);
   VitalWireDelay (B1_ipd, B1, tipd_B1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((B0_ipd) AND (A0_ipd) AND (A1_ipd)) OR ((B1_ipd) AND (A1_ipd)) OR
         ((B0_ipd) AND (A0_ipd) AND (B1_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B1_ipd'last_event, tpd_B1_Y, TRUE),
                 1 => (B0_ipd'last_event, tpd_B0_Y, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_Y, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CY2A_VITAL of CY2A is
   for VITAL_ACT
   end for;
end CFG_CY2A_VITAL;


----- CELL CY2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CY2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CY2B : entity is TRUE;
end CY2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of CY2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B0_ipd, B0, tipd_B0);
   VitalWireDelay (B1_ipd, B1, tipd_B1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((A1_ipd) AND ((B0_ipd) OR (A0_ipd))) OR ((B1_ipd) AND (A1_ipd)) OR
         ((B1_ipd) AND ((B0_ipd) OR (A0_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B1_ipd'last_event, tpd_B1_Y, TRUE),
                 1 => (B0_ipd'last_event, tpd_B0_Y, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_Y, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CY2B_VITAL of CY2B is
   for VITAL_ACT
   end for;
end CFG_CY2B_VITAL;










----- CELL DECETH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity DECETH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF DECETH : ENTITY IS TRUE;
	--
end DECETH;

ARCHITECTURE VITAL_ACT OF DECETH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  DECETH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  DECETH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  DECETH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 5);
		--VARIABLE  PrevData_DECETH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_DECETH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : DECETH_TAB Declaration
		CONSTANT  DECETH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
                --Vio, Clr, Clk,   d,   e, prev, next 
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_ODE_CLK or 
				SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : DECETH_TAB
		VitalStateTable (
				StateTable         => DECETH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => DFE3C_Result,
				PreviousDataIn     => PrevData_DFE3C
		);	--End VitalStateTable
		DFE3CStateReg(0)          := DFE3C_Result(2);
		IQ(0)                     := DFE3C_Result(1);
		--
		--Implement Functionality for State Table : DECETH_TAB
		VitalStateTable (
				StateTable         => DECETH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & PAD_ipd & IDE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_ipd, IDE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => DECETH_TAB_Result,
				PreviousDataIn     => PrevData_DECETH_TAB
		);	--End VitalStateTable
		DECETH_TABStateReg(0)     := DECETH_TAB_Result(2);
		Q_zd                      := DECETH_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;


		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_DECETH_VITAL of DECETH is
   for VITAL_ACT
   end for;
end CFG_DECETH_VITAL;
----- CELL DECETL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity DECETL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Removal time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF DECETL : ENTITY IS TRUE;
	--
end DECETL;

ARCHITECTURE VITAL_ACT OF DECETL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  DECETL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  DECETL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  DECETL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 5);
		--VARIABLE  PrevData_DECETL_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_DECETL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : DECETL_TAB Declaration
		CONSTANT  DECETL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_ODE_CLK or 
				SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : DECETL_TAB
		VitalStateTable (
				StateTable         => DECETL_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => DFE3C_Result,
				PreviousDataIn     => PrevData_DFE3C
		);	--End VitalStateTable
		DFE3CStateReg(0)          := DFE3C_Result(2);
		IQ(0)                     := DFE3C_Result(1);
		--
		--Implement Functionality for State Table : DECETL_TAB
		VitalStateTable (
				StateTable         => DECETL_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & PAD_ipd & IDE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_ipd, IDE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => DECETL_TAB_Result,
				PreviousDataIn     => PrevData_DECETL_TAB
		);	--End VitalStateTable
		DECETL_TABStateReg(0)     := DECETL_TAB_Result(2);
		Q_zd                      := DECETL_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_DECETL_VITAL of DECETL is
   for VITAL_ACT
   end for;
end CFG_DECETL_VITAL;
----- CELL DEPETH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity DEPETH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF DEPETH : ENTITY IS TRUE;
	--
end DEPETH;

ARCHITECTURE VITAL_ACT OF DEPETH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  DEPETH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  DEPETH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  DEPETH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 5);
		--VARIABLE  PrevData_DEPETH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_DEPETH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : DEPETH_TAB Declaration
		CONSTANT  DEPETH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
--          Violation, IOPCL, CLK, D, ODE
		( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_ODE_CLK or 
				SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : DEPETH_TAB
		VitalStateTable (
				StateTable         => DEPETH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => DFE3C_Result,
				PreviousDataIn     => PrevData_DFE3C
		);	--End VitalStateTable
		DFE3CStateReg(0)          := DFE3C_Result(2);
		IQ(0)                     := DFE3C_Result(1);
		--
		--Implement Functionality for State Table : DEPETH_TAB
		VitalStateTable (
				StateTable         => DEPETH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & PAD_ipd & IDE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_ipd, IDE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => DEPETH_TAB_Result,
				PreviousDataIn     => PrevData_DEPETH_TAB
		);	--End VitalStateTable
		DEPETH_TABStateReg(0)     := DEPETH_TAB_Result(2);
		Q_zd                      := DEPETH_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_DEPETH_VITAL of DEPETH is
   for VITAL_ACT
   end for;
end CFG_DEPETH_VITAL;
----- CELL DEPETL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity DEPETL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_Q          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Q
		tpd_CLK_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Q
		tpd_PAD_Q            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Q
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IDE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IDE
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between PAD and CLK
		tsetup_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between IDE and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_PAD_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between PAD and CLK
		thold_IDE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IDE and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IDE                 : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Q                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF DEPETL : ENTITY IS TRUE;
	--
end DEPETL;

ARCHITECTURE VITAL_ACT OF DEPETL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IDE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IDE_ipd,
				InSig              => IDE,
				twire              => tipd_IDE
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IDE_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  PAD_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  IDE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Q_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_PAD_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_IDE_CLK              : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  DFE3CStateReg             : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  IQ                        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  DEPETL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  DFE3C_Result              : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		VARIABLE  DEPETL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  DEPETL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 5);
		--VARIABLE  PrevData_DEPETL_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_DFE3C            : STD_LOGIC_VECTOR(0 TO 4);
		VARIABLE  PrevData_DEPETL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Q_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		VARIABLE  IDE_delayed               : STD_ULOGIC;
		VARIABLE  PAD_delayed               : STD_ULOGIC;
		--
		-- State Table : DEPETL_TAB Declaration
		CONSTANT  DEPETL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
--          Violation, IOPCL, CLK, D, ODE
		( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : PAD
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_PAD_CLK,
				TimingData         => PAD_CLK_TimingDataSH,
				TestSignal         => PAD_ipd,
				TestSignalName     => "PAD",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_PAD_CLK_noedge_posedge,
				SetupLow           => tsetup_PAD_CLK_noedge_posedge,
				HoldHigh           => thold_PAD_CLK_noedge_posedge,
				HoldLow            => thold_PAD_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR IDE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : IDE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_IDE_CLK,
				TimingData         => IDE_CLK_TimingDataSH,
				TestSignal         => IDE_ipd,
				TestSignalName     => "IDE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_IDE_CLK_noedge_posedge,
				SetupLow           => tsetup_IDE_CLK_noedge_posedge,
				HoldHigh           => thold_IDE_CLK_noedge_posedge,
				HoldLow            => thold_IDE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_IDE_CLK or SHVF_ODE_CLK or 
				SHVF_PAD_CLK ;
		--
		--Implement Functionality for State Table : DEPETL_TAB
		VitalStateTable (
				StateTable         => DEPETL_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => DFE3C_Result,
				PreviousDataIn     => PrevData_DFE3C
		);	--End VitalStateTable
		DFE3CStateReg(0)          := DFE3C_Result(2);
		IQ(0)                     := DFE3C_Result(1);
		--
		--Implement Functionality for State Table : DEPETL_TAB
		VitalStateTable (
				StateTable         => DEPETL_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & PAD_ipd & IDE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_ipd, IDE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, PAD_delayed, IDE_delayed),
				NumStates          => 1,
				Result             => DEPETL_TAB_Result,
				PreviousDataIn     => PrevData_DEPETL_TAB
		);	--End VitalStateTable
		DEPETL_TABStateReg(0)     := DEPETL_TAB_Result(2);
		Q_zd                      := DEPETL_TAB_Result(1);
		--
		PAD_zd := VitalBUFIF0 (data => IQ(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;
		IDE_delayed := IDE_ipd;
		PAD_delayed := PAD_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Q,
				OutSignalName      => "Q",
				OutTemp            => Q_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Q,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Q,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Q,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Q_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_DEPETL_VITAL of DEPETL is
   for VITAL_ACT
   end for;
end CFG_DEPETL_VITAL;
----- CELL DF1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1 : entity is TRUE;
end DF1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1_VITAL of DF1 is
   for VITAL_ACT
   end for;
end CFG_DF1_VITAL;


----- CELL DF1_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1_CC : entity is TRUE;
end DF1_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1_CC_VITAL of DF1_CC is
   for VITAL_ACT
   end for;
end CFG_DF1_CC_VITAL;


----- CELL DF1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1A : entity is TRUE;
end DF1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1A_VITAL of DF1A is
   for VITAL_ACT
   end for;
end CFG_DF1A_VITAL;


----- CELL DF1A_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1A_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1A_CC : entity is TRUE;
end DF1A_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1A_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1A_CC_VITAL of DF1A_CC is
   for VITAL_ACT
   end for;
end CFG_DF1A_CC_VITAL;


----- CELL DF1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1B : entity is TRUE;
end DF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1B_VITAL of DF1B is
   for VITAL_ACT
   end for;
end CFG_DF1B_VITAL;


----- CELL DF1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1B_CC : entity is TRUE;
end DF1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1B_CC_VITAL of DF1B_CC is
   for VITAL_ACT
   end for;
end CFG_DF1B_CC_VITAL;


----- CELL DF1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1C : entity is TRUE;
end DF1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1C_VITAL of DF1C is
   for VITAL_ACT
   end for;
end CFG_DF1C_VITAL;


----- CELL DF1C_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1C_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1C_CC : entity is TRUE;
end DF1C_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DF1C_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1C_CC_VITAL of DF1C_CC is
   for VITAL_ACT
   end for;
end CFG_DF1C_CC_VITAL;


----- CELL DFC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1 : entity is TRUE;
end DFC1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)


   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1_VITAL of DFC1 is
   for VITAL_ACT
   end for;
end CFG_DFC1_VITAL;


----- CELL DFC1_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1_CC : entity is TRUE;
end DFC1_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1_CC_VITAL of DFC1_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1_CC_VITAL;


----- CELL DFC1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1A : entity is TRUE;
end DFC1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1A_VITAL of DFC1A is
   for VITAL_ACT
   end for;
end CFG_DFC1A_VITAL;


----- CELL DFC1A_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1A_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1A_CC : entity is TRUE;
end DFC1A_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1A_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1A_CC_VITAL of DFC1A_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1A_CC_VITAL;


----- CELL DFC1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1B : entity is TRUE;
end DFC1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1B_VITAL of DFC1B is
   for VITAL_ACT
   end for;
end CFG_DFC1B_VITAL;


----- CELL DFC1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1B_CC : entity is TRUE;
end DFC1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_CC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_CC_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1B_CC_VITAL of DFC1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1B_CC_VITAL;


----- CELL DFC1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1D : entity is TRUE;
end DFC1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1D_VITAL of DFC1D is
   for VITAL_ACT
   end for;
end CFG_DFC1D_VITAL;


----- CELL DFC1D_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1D_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1D_CC : entity is TRUE;
end DFC1D_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1D_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1D_CC_VITAL of DFC1D_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1D_CC_VITAL;


----- CELL DFC1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1E : entity is TRUE;
end DFC1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1E_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  H,  x,  L ),
    ( L,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( x,  L,  x,  x,  x,  H ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  U,  x,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFC1E_QN_tab,
        DataIn => (
               CLK_delayed, CLR_ipd, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1E_VITAL of DFC1E is
   for VITAL_ACT
   end for;
end CFG_DFC1E_VITAL;


----- CELL DFC1G -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1G is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1G : entity is TRUE;
end DFC1G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1G is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1E_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  H,  x,  L ),
    ( L,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( x,  L,  x,  x,  x,  H ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  U,  x,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFC1E_QN_tab,
        DataIn => (
               CLK_ipd, CLR_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1G_VITAL of DFC1G is
   for VITAL_ACT
   end for;
end CFG_DFC1G_VITAL;


----- CELL DFE -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE : entity is TRUE;
end DFE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE_VITAL of DFE is
   for VITAL_ACT
   end for;
end CFG_DFE_VITAL;


----- CELL DFE_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE_CC : entity is TRUE;
end DFE_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE_CC_VITAL of DFE_CC is
   for VITAL_ACT
   end for;
end CFG_DFE_CC_VITAL;


----- CELL DFE1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1B : entity is TRUE;
end DFE1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1B_VITAL of DFE1B is
   for VITAL_ACT
   end for;
end CFG_DFE1B_VITAL;


----- CELL DFE1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1B_CC : entity is TRUE;
end DFE1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)


   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1B_CC_VITAL of DFE1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFE1B_CC_VITAL;


----- CELL DFE1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1C : entity is TRUE;
end DFE1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0' ,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1C_VITAL of DFE1C is
   for VITAL_ACT
   end for;
end CFG_DFE1C_VITAL;


----- CELL DFE1C_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1C_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1C_CC : entity is TRUE;
end DFE1C_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1C_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0' ,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1C_CC_VITAL of DFE1C_CC is
   for VITAL_ACT
   end for;
end CFG_DFE1C_CC_VITAL;


----- CELL DFE3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3A : entity is TRUE;
end DFE3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  H,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( CLR_ipd ) AND ( E_ipd )) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3A_VITAL of DFE3A is
   for VITAL_ACT
   end for;
end CFG_DFE3A_VITAL;


----- CELL DFE3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3B : entity is TRUE;
end DFE3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  H,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( CLR_ipd ) AND ( E_ipd )) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3B_VITAL of DFE3B is
   for VITAL_ACT
   end for;
end CFG_DFE3B_VITAL;


----- CELL DFE3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3C : entity is TRUE;
end DFE3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3C_VITAL of DFE3C is
   for VITAL_ACT
   end for;
end CFG_DFE3C_VITAL;


----- CELL DFE3D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3D : entity is TRUE;
end DFE3D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3D_VITAL of DFE3D is
   for VITAL_ACT
   end for;
end CFG_DFE3D_VITAL;


----- CELL DFEA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEA : entity is TRUE;
end DFEA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFEA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFEA_VITAL of DFEA is
   for VITAL_ACT
   end for;
end CFG_DFEA_VITAL;


----- CELL DFEA_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEA_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEA_CC : entity is TRUE;
end DFEA_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFEA_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFEA_CC_VITAL of DFEA_CC is
   for VITAL_ACT
   end for;
end CFG_DFEA_CC_VITAL;


----- CELL DFM -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM : entity is TRUE;
end DFM;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM_VITAL of DFM is
   for VITAL_ACT
   end for;
end CFG_DFM_VITAL;


----- CELL DFM_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM_CC : entity is TRUE;
end DFM_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM_CC_VITAL of DFM_CC is
   for VITAL_ACT
   end for;
end CFG_DFM_CC_VITAL;


----- CELL DFM1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1B : entity is TRUE;
end DFM1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_QN_tab,
        DataIn => (
               CLK_delayed, S_delayed, B_delayed, A_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1B_VITAL of DFM1B is
   for VITAL_ACT
   end for;
end CFG_DFM1B_VITAL;


----- CELL DFM1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1B_CC : entity is TRUE;
end DFM1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_CC_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_CC_QN_tab,
        DataIn => (
               CLK_delayed, S_delayed, B_delayed, A_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1B_CC_VITAL of DFM1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFM1B_CC_VITAL;


----- CELL DFM1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1C : entity is TRUE;
end DFM1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_QN_tab,
        DataIn => (
               CLK_ipd, S_delayed, B_delayed, A_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1C_VITAL of DFM1C is
   for VITAL_ACT
   end for;
end CFG_DFM1C_VITAL;


----- CELL DFM1C_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1C_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1C_CC : entity is TRUE;
end DFM1C_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1C_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_QN_tab,
        DataIn => (
               CLK_ipd, S_delayed, B_delayed, A_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1C_CC_VITAL of DFM1C_CC is
   for VITAL_ACT
   end for;
end CFG_DFM1C_CC_VITAL;


----- CELL DFM3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM3 : entity is TRUE;
end DFM3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLR or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM3_VITAL of DFM3 is
   for VITAL_ACT
   end for;
end CFG_DFM3_VITAL;


----- CELL DFM3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM3B : entity is TRUE;
end DFM3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM3B_VITAL of DFM3B is
   for VITAL_ACT
   end for;
end CFG_DFM3B_VITAL;


----- CELL DFM3E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM3E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM3E : entity is TRUE;
end DFM3E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM3E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM3E_VITAL of DFM3E is
   for VITAL_ACT
   end for;
end CFG_DFM3E_VITAL;


----- CELL DFM4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM4C : entity is TRUE;
end DFM4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM4C_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  H,  H,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM4C_QN_tab,
        DataIn => (
               PRE_ipd, CLK_delayed, S_delayed, B_delayed, A_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM4C_VITAL of DFM4C is
   for VITAL_ACT
   end for;
end CFG_DFM4C_VITAL;


----- CELL DFM4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM4D : entity is TRUE;
end DFM4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM4C_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  H,  H,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Pviol_PRE or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM4C_QN_tab,
        DataIn => (
               PRE_ipd, CLK_ipd, S_delayed, B_delayed, A_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM4D_VITAL of DFM4D is
   for VITAL_ACT
   end for;
end CFG_DFM4D_VITAL;


----- CELL DFM6A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM6A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM6A : entity is TRUE;
end DFM6A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM6A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S1_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM6A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_posedge,
          TimingData              => Tmkr_D0_CLK_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_posedge,
          SetupLow                => tsetup_D0_CLK_noedge_posedge,
          HoldHigh                => thold_D0_CLK_noedge_posedge,
          HoldLow                 => thold_D0_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_posedge,
          TimingData              => Tmkr_D1_CLK_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_posedge,
          SetupLow                => tsetup_D1_CLK_noedge_posedge,
          HoldHigh                => thold_D1_CLK_noedge_posedge,
          HoldLow                 => thold_D1_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_posedge,
          TimingData              => Tmkr_D2_CLK_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_posedge,
          SetupLow                => tsetup_D2_CLK_noedge_posedge,
          HoldHigh                => thold_D2_CLK_noedge_posedge,
          HoldLow                 => thold_D2_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_posedge,
          TimingData              => Tmkr_D3_CLK_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_posedge,
          SetupLow                => tsetup_D3_CLK_noedge_posedge,
          HoldHigh                => thold_D3_CLK_noedge_posedge,
          HoldLow                 => thold_D3_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_posedge,
          TimingData              => Tmkr_S0_CLK_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_posedge,
          SetupLow                => tsetup_S0_CLK_noedge_posedge,
          HoldHigh                => thold_S0_CLK_noedge_posedge,
          HoldLow                 => thold_S0_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_CLK_posedge,
          TimingData              => Tmkr_S1_CLK_posedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_CLK_noedge_posedge,
          SetupLow                => tsetup_S1_CLK_noedge_posedge,
          HoldHigh                => thold_S1_CLK_noedge_posedge,
          HoldLow                 => thold_S1_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_posedge or Tviol_D3_CLK_posedge or Tviol_S1_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_D1_CLK_posedge or Tviol_D2_CLK_posedge or Tviol_S0_CLK_posedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM6A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S1_delayed, S0_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S1_delayed := S1_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM6A_VITAL of DFM6A is
   for VITAL_ACT
   end for;
end CFG_DFM6A_VITAL;


----- CELL DFM6B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM6B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM6B : entity is TRUE;
end DFM6B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM6B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S1_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM6A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_negedge,
          TimingData              => Tmkr_D0_CLK_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_negedge,
          SetupLow                => tsetup_D0_CLK_noedge_negedge,
          HoldHigh                => thold_D0_CLK_noedge_negedge,
          HoldLow                 => thold_D0_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_negedge,
          TimingData              => Tmkr_D1_CLK_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_negedge,
          SetupLow                => tsetup_D1_CLK_noedge_negedge,
          HoldHigh                => thold_D1_CLK_noedge_negedge,
          HoldLow                 => thold_D1_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_negedge,
          TimingData              => Tmkr_D2_CLK_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_negedge,
          SetupLow                => tsetup_D2_CLK_noedge_negedge,
          HoldHigh                => thold_D2_CLK_noedge_negedge,
          HoldLow                 => thold_D2_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_negedge,
          TimingData              => Tmkr_D3_CLK_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_negedge,
          SetupLow                => tsetup_D3_CLK_noedge_negedge,
          HoldHigh                => thold_D3_CLK_noedge_negedge,
          HoldLow                 => thold_D3_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_negedge,
          TimingData              => Tmkr_S0_CLK_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_negedge,
          SetupLow                => tsetup_S0_CLK_noedge_negedge,
          HoldHigh                => thold_S0_CLK_noedge_negedge,
          HoldLow                 => thold_S0_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_CLK_negedge,
          TimingData              => Tmkr_S1_CLK_negedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_CLK_noedge_negedge,
          SetupLow                => tsetup_S1_CLK_noedge_negedge,
          HoldHigh                => thold_S1_CLK_noedge_negedge,
          HoldLow                 => thold_S1_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_negedge or Tviol_D1_CLK_negedge or Tviol_D2_CLK_negedge or Tviol_S0_CLK_negedge or Tviol_D3_CLK_negedge or Tviol_S1_CLK_negedge or Pviol_CLR or Tviol_CLR_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM6A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S1_delayed, S0_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S1_delayed := S1_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM6B_VITAL of DFM6B is
   for VITAL_ACT
   end for;
end CFG_DFM6B_VITAL;


----- CELL DFM7A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM7A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM7A : entity is TRUE;
end DFM7A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM7A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 9);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S10_delayed : STD_ULOGIC := 'X';
   VARIABLE S11_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM7A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_posedge,
          TimingData              => Tmkr_D0_CLK_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_posedge,
          SetupLow                => tsetup_D0_CLK_noedge_posedge,
          HoldHigh                => thold_D0_CLK_noedge_posedge,
          HoldLow                 => thold_D0_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_posedge,
          TimingData              => Tmkr_D1_CLK_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_posedge,
          SetupLow                => tsetup_D1_CLK_noedge_posedge,
          HoldHigh                => thold_D1_CLK_noedge_posedge,
          HoldLow                 => thold_D1_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_posedge,
          TimingData              => Tmkr_D2_CLK_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_posedge,
          SetupLow                => tsetup_D2_CLK_noedge_posedge,
          HoldHigh                => thold_D2_CLK_noedge_posedge,
          HoldLow                 => thold_D2_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_posedge,
          TimingData              => Tmkr_D3_CLK_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_posedge,
          SetupLow                => tsetup_D3_CLK_noedge_posedge,
          HoldHigh                => thold_D3_CLK_noedge_posedge,
          HoldLow                 => thold_D3_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_posedge,
          TimingData              => Tmkr_S0_CLK_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_posedge,
          SetupLow                => tsetup_S0_CLK_noedge_posedge,
          HoldHigh                => thold_S0_CLK_noedge_posedge,
          HoldLow                 => thold_S0_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_CLK_posedge,
          TimingData              => Tmkr_S10_CLK_posedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_CLK_noedge_posedge,
          SetupLow                => tsetup_S10_CLK_noedge_posedge,
          HoldHigh                => thold_S10_CLK_noedge_posedge,
          HoldLow                 => thold_S10_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_CLK_posedge,
          TimingData              => Tmkr_S11_CLK_posedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_CLK_noedge_posedge,
          SetupLow                => tsetup_S11_CLK_noedge_posedge,
          HoldHigh                => thold_S11_CLK_noedge_posedge,
          HoldLow                 => thold_S11_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_posedge or Tviol_D3_CLK_posedge or Tviol_S11_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_D1_CLK_posedge or Tviol_D2_CLK_posedge or Tviol_S0_CLK_posedge or Pviol_CLR or Tviol_S10_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM7A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S11_delayed, S10_delayed, S0_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S10_delayed := S10_ipd;
      S11_delayed := S11_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM7A_VITAL of DFM7A is
   for VITAL_ACT
   end for;
end CFG_DFM7A_VITAL;


----- CELL DFM7B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM7B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM7B : entity is TRUE;
end DFM7B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM7B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 9);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S10_delayed : STD_ULOGIC := 'X';
   VARIABLE S11_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM7A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_negedge,
          TimingData              => Tmkr_D0_CLK_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_negedge,
          SetupLow                => tsetup_D0_CLK_noedge_negedge,
          HoldHigh                => thold_D0_CLK_noedge_negedge,
          HoldLow                 => thold_D0_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_negedge,
          TimingData              => Tmkr_D1_CLK_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_negedge,
          SetupLow                => tsetup_D1_CLK_noedge_negedge,
          HoldHigh                => thold_D1_CLK_noedge_negedge,
          HoldLow                 => thold_D1_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_negedge,
          TimingData              => Tmkr_D2_CLK_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_negedge,
          SetupLow                => tsetup_D2_CLK_noedge_negedge,
          HoldHigh                => thold_D2_CLK_noedge_negedge,
          HoldLow                 => thold_D2_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_negedge,
          TimingData              => Tmkr_D3_CLK_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_negedge,
          SetupLow                => tsetup_D3_CLK_noedge_negedge,
          HoldHigh                => thold_D3_CLK_noedge_negedge,
          HoldLow                 => thold_D3_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_negedge,
          TimingData              => Tmkr_S0_CLK_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_negedge,
          SetupLow                => tsetup_S0_CLK_noedge_negedge,
          HoldHigh                => thold_S0_CLK_noedge_negedge,
          HoldLow                 => thold_S0_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_CLK_negedge,
          TimingData              => Tmkr_S10_CLK_negedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_CLK_noedge_negedge,
          SetupLow                => tsetup_S10_CLK_noedge_negedge,
          HoldHigh                => thold_S10_CLK_noedge_negedge,
          HoldLow                 => thold_S10_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_CLK_negedge,
          TimingData              => Tmkr_S11_CLK_negedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_CLK_noedge_negedge,
          SetupLow                => tsetup_S11_CLK_noedge_negedge,
          HoldHigh                => thold_S11_CLK_noedge_negedge,
          HoldLow                 => thold_S11_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_negedge or Tviol_D1_CLK_negedge or Tviol_D2_CLK_negedge or Tviol_S0_CLK_negedge or Tviol_S10_CLK_negedge or Tviol_D3_CLK_negedge or Pviol_CLR or Tviol_S11_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM7A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S11_delayed, S10_delayed, S0_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S10_delayed := S10_ipd;
      S11_delayed := S11_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM7B_VITAL of DFM7B is
   for VITAL_ACT
   end for;
end CFG_DFM7B_VITAL;


----- CELL DFM8A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM8A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S00_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S00_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S01_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S01_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S00                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S01                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM8A : entity is TRUE;
end DFM8A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM8A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S00_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S01_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S00_ipd, S00, tipd_S00);
   VitalWireDelay (S01_ipd, S01, tipd_S01);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S00_ipd, S01_ipd, S10_ipd, S11_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S00_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S00_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S01_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S01_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 10);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S00_delayed : STD_ULOGIC := 'X';
   VARIABLE S01_delayed : STD_ULOGIC := 'X';
   VARIABLE S10_delayed : STD_ULOGIC := 'X';
   VARIABLE S11_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM8A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_posedge,
          TimingData              => Tmkr_D0_CLK_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_posedge,
          SetupLow                => tsetup_D0_CLK_noedge_posedge,
          HoldHigh                => thold_D0_CLK_noedge_posedge,
          HoldLow                 => thold_D0_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_posedge,
          TimingData              => Tmkr_D1_CLK_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_posedge,
          SetupLow                => tsetup_D1_CLK_noedge_posedge,
          HoldHigh                => thold_D1_CLK_noedge_posedge,
          HoldLow                 => thold_D1_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd ))
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_posedge,
          TimingData              => Tmkr_D2_CLK_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_posedge,
          SetupLow                => tsetup_D2_CLK_noedge_posedge,
          HoldHigh                => thold_D2_CLK_noedge_posedge,
          HoldLow                 => thold_D2_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_posedge,
          TimingData              => Tmkr_D3_CLK_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_posedge,
          SetupLow                => tsetup_D3_CLK_noedge_posedge,
          HoldHigh                => thold_D3_CLK_noedge_posedge,
          HoldLow                 => thold_D3_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd ))
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S00_CLK_posedge,
          TimingData              => Tmkr_S00_CLK_posedge,
          TestSignal              => S00_ipd,
          TestSignalName          => "S00",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S00_CLK_noedge_posedge,
          SetupLow                => tsetup_S00_CLK_noedge_posedge,
          HoldHigh                => thold_S00_CLK_noedge_posedge,
          HoldLow                 => thold_S00_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S01_CLK_posedge,
          TimingData              => Tmkr_S01_CLK_posedge,
          TestSignal              => S01_ipd,
          TestSignalName          => "S01",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S01_CLK_noedge_posedge,
          SetupLow                => tsetup_S01_CLK_noedge_posedge,
          HoldHigh                => thold_S01_CLK_noedge_posedge,
          HoldLow                 => thold_S01_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_CLK_posedge,
          TimingData              => Tmkr_S10_CLK_posedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_CLK_noedge_posedge,
          SetupLow                => tsetup_S10_CLK_noedge_posedge,
          HoldHigh                => thold_S10_CLK_noedge_posedge,
          HoldLow                 => thold_S10_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_CLK_posedge,
          TimingData              => Tmkr_S11_CLK_posedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_CLK_noedge_posedge,
          SetupLow                => tsetup_S11_CLK_noedge_posedge,
          HoldHigh                => thold_S11_CLK_noedge_posedge,
          HoldLow                 => thold_S11_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_posedge or Tviol_D3_CLK_posedge or Tviol_S00_CLK_posedge or Tviol_S11_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_D1_CLK_posedge or Tviol_D2_CLK_posedge or Tviol_S01_CLK_posedge or Tviol_S10_CLK_posedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM8A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D2_delayed, D3_delayed, D0_delayed, D1_delayed, S11_delayed, S10_delayed, S01_delayed, S00_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S00_delayed := S00_ipd;
      S01_delayed := S01_ipd;
      S10_delayed := S10_ipd;
      S11_delayed := S11_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM8A_VITAL of DFM8A is
   for VITAL_ACT
   end for;
end CFG_DFM8A_VITAL;


----- CELL DFM8B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM8B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S00_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S00_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S01_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S01_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM8B : entity is TRUE;
end DFM8B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM8B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S00_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S01_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S00_ipd, S00, tipd_S00);
   VitalWireDelay (S01_ipd, S01, tipd_S01);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S00_ipd, S01_ipd, S10_ipd, S11_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S00_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S00_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S01_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S01_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 10);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S00_delayed : STD_ULOGIC := 'X';
   VARIABLE S01_delayed : STD_ULOGIC := 'X';
   VARIABLE S10_delayed : STD_ULOGIC := 'X';
   VARIABLE S11_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM8A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_negedge,
          TimingData              => Tmkr_D0_CLK_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_negedge,
          SetupLow                => tsetup_D0_CLK_noedge_negedge,
          HoldHigh                => thold_D0_CLK_noedge_negedge,
          HoldLow                 => thold_D0_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd ) 
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_negedge,
          TimingData              => Tmkr_D1_CLK_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_negedge,
          SetupLow                => tsetup_D1_CLK_noedge_negedge,
          HoldHigh                => thold_D1_CLK_noedge_negedge,
          HoldLow                 => thold_D1_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd )) 
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_negedge,
          TimingData              => Tmkr_D2_CLK_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_negedge,
          SetupLow                => tsetup_D2_CLK_noedge_negedge,
          HoldHigh                => thold_D2_CLK_noedge_negedge,
          HoldLow                 => thold_D2_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd ) 
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_negedge,
          TimingData              => Tmkr_D3_CLK_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_negedge,
          SetupLow                => tsetup_D3_CLK_noedge_negedge,
          HoldHigh                => thold_D3_CLK_noedge_negedge,
          HoldLow                 => thold_D3_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd )) 
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S00_CLK_negedge,
          TimingData              => Tmkr_S00_CLK_negedge,
          TestSignal              => S00_ipd,
          TestSignalName          => "S00",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S00_CLK_noedge_negedge,
          SetupLow                => tsetup_S00_CLK_noedge_negedge,
          HoldHigh                => thold_S00_CLK_noedge_negedge,
          HoldLow                 => thold_S00_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S01_CLK_negedge,
          TimingData              => Tmkr_S01_CLK_negedge,
          TestSignal              => S01_ipd,
          TestSignalName          => "S01",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S01_CLK_noedge_negedge,
          SetupLow                => tsetup_S01_CLK_noedge_negedge,
          HoldHigh                => thold_S01_CLK_noedge_negedge,
          HoldLow                 => thold_S01_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_CLK_negedge,
          TimingData              => Tmkr_S10_CLK_negedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_CLK_noedge_negedge,
          SetupLow                => tsetup_S10_CLK_noedge_negedge,
          HoldHigh                => thold_S10_CLK_noedge_negedge,
          HoldLow                 => thold_S10_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_CLK_negedge,
          TimingData              => Tmkr_S11_CLK_negedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_CLK_noedge_negedge,
          SetupLow                => tsetup_S11_CLK_noedge_negedge,
          HoldHigh                => thold_S11_CLK_noedge_negedge,
          HoldLow                 => thold_S11_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_negedge or Tviol_D1_CLK_negedge or Tviol_D2_CLK_negedge or Tviol_S01_CLK_negedge or Tviol_S10_CLK_negedge or Tviol_D3_CLK_negedge or Pviol_CLR or Tviol_S00_CLK_negedge or Tviol_CLR_CLK_negedge or Tviol_S11_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM8A_Q_tab,
        DataIn => (
               CLR_ipd, ( NOT CLK_delayed ), D2_delayed, D3_delayed, D0_delayed, D1_delayed, S11_delayed, S10_delayed, S01_delayed, S00_delayed, (NOT CLK_ipd )));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S00_delayed := S00_ipd;
      S01_delayed := S01_ipd;
      S10_delayed := S10_ipd;
      S11_delayed := S11_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM8B_VITAL of DFM8B is
   for VITAL_ACT
   end for;
end CFG_DFM8B_VITAL;


----- CELL DFMA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFMA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFMA : entity is TRUE;
end DFMA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFMA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFMA_VITAL of DFMA is
   for VITAL_ACT
   end for;
end CFG_DFMA_VITAL;


----- CELL DFMA_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFMA_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFMA_CC : entity is TRUE;
end DFMA_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFMA_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFMA_CC_VITAL of DFMA_CC is
   for VITAL_ACT
   end for;
end CFG_DFMA_CC_VITAL;


----- CELL DFMB -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFMB is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFMB : entity is TRUE;
end DFMB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFMB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLR or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFMB_VITAL of DFMB is
   for VITAL_ACT
   end for;
end CFG_DFMB_VITAL;


----- CELL DFME1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFME1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFME1A : entity is TRUE;
end DFME1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFME1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H,  L,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  H,  x,  H,  L,  H,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR (NOT S_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_E_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFME1A_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, B_delayed, A_delayed, S_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFME1A_VITAL of DFME1A is
   for VITAL_ACT
   end for;
end CFG_DFME1A_VITAL;


----- CELL DFP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1 : entity is TRUE;
end DFP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1_VITAL of DFP1 is
   for VITAL_ACT
   end for;
end CFG_DFP1_VITAL;


----- CELL DFP1_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1_CC : entity is TRUE;
end DFP1_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_CC_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_CC_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1_CC_VITAL of DFP1_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1_CC_VITAL;


----- CELL DFP1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1A : entity is TRUE;
end DFP1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1A_VITAL of DFP1A is
   for VITAL_ACT
   end for;
end CFG_DFP1A_VITAL;


----- CELL DFP1A_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1A_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1A_CC : entity is TRUE;
end DFP1A_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1A_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1A_CC_VITAL of DFP1A_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1A_CC_VITAL;


----- CELL DFP1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1B : entity is TRUE;
end DFP1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1B_VITAL of DFP1B is
   for VITAL_ACT
   end for;
end CFG_DFP1B_VITAL;


----- CELL DFP1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1B_CC : entity is TRUE;
end DFP1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_CC_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_CC_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1B_CC_VITAL of DFP1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1B_CC_VITAL;


----- CELL DFP1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1C : entity is TRUE;
end DFP1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1C_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  L,  x,  H ),
    ( L,  H,  H,  x,  x,  L ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1C_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd, PRE_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1C_VITAL of DFP1C is
   for VITAL_ACT
   end for;
end CFG_DFP1C_VITAL;


----- CELL DFP1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1D : entity is TRUE;
end DFP1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1D_VITAL of DFP1D is
   for VITAL_ACT
   end for;
end CFG_DFP1D_VITAL;


----- CELL DFP1D_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1D_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1D_CC : entity is TRUE;
end DFP1D_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1D_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1D_CC_VITAL of DFP1D_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1D_CC_VITAL;


----- CELL DFP1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1E : entity is TRUE;
end DFP1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1E_QN_tab,
        DataIn => (
               PRE_ipd, CLK_delayed, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1E_VITAL of DFP1E is
   for VITAL_ACT
   end for;
end CFG_DFP1E_VITAL;


----- CELL DFP1F -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1F is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1F : entity is TRUE;
end DFP1F;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1F is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1C_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  L,  x,  H ),
    ( L,  H,  H,  x,  x,  L ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1C_QN_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed, PRE_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1F_VITAL of DFP1F is
   for VITAL_ACT
   end for;
end CFG_DFP1F_VITAL;


----- CELL DFP1G -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1G is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1G : entity is TRUE;
end DFP1G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1G is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1E_QN_tab,
        DataIn => (
               PRE_ipd, CLK_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1G_VITAL of DFP1G is
   for VITAL_ACT
   end for;
end CFG_DFP1G_VITAL;


----- CELL DFPC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPC : entity is TRUE;
end DFPC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_PRE or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPC_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPC_VITAL of DFPC is
   for VITAL_ACT
   end for;
end CFG_DFPC_VITAL;


----- CELL DFPC_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPC_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPC_CC : entity is TRUE;
end DFPC_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPC_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPC_CC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_PRE or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPC_CC_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPC_CC_VITAL of DFPC_CC is
   for VITAL_ACT
   end for;
end CFG_DFPC_CC_VITAL;


----- CELL DFPCA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPCA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPCA : entity is TRUE;
end DFPCA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPCA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPCA_tab : VitalStateTableType := (
    ( L,  x,  x,  H,  x,  x,  U ),
    ( L,  x,  x,  L,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPCA_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPCA_VITAL of DFPCA is
   for VITAL_ACT
   end for;
end CFG_DFPCA_VITAL;


----- CELL DFPCA_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPCA_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPCA_CC : entity is TRUE;
end DFPCA_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPCA_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPCA_CC_tab : VitalStateTableType := (
    ( L,  x,  x,  H,  x,  x,  U ),
    ( L,  x,  x,  L,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPCA_CC_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPCA_CC_VITAL of DFPCA_CC is
   for VITAL_ACT
   end for;
end CFG_DFPCA_CC_VITAL;


----- CELL DL1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1 : entity is TRUE;
end DL1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DL1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1_Q_tab,
        DataIn => (
               D_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1_VITAL of DL1 is
   for VITAL_ACT
   end for;
end CFG_DL1_VITAL;


----- CELL DL1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1A : entity is TRUE;
end DL1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DL1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL1A_QN_tab,
        DataIn => (
               D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1A_VITAL of DL1A is
   for VITAL_ACT
   end for;
end CFG_DL1A_VITAL;


----- CELL DL1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1B : entity is TRUE;
end DL1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DL1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1B_Q_tab,
        DataIn => (
               G_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1B_VITAL of DL1B is
   for VITAL_ACT
   end for;
end CFG_DL1B_VITAL;


----- CELL DL1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1C : entity is TRUE;
end DL1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DL1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL1C_QN_tab,
        DataIn => (
               G_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1C_VITAL of DL1C is
   for VITAL_ACT
   end for;
end CFG_DL1C_VITAL;


----- CELL DL2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2A : entity is TRUE;
end DL2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  L,  x,  S ),
    ( H,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ),
    ( H,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL2A_Q_tab,
        DataIn => (
               CLR_ipd, D_ipd, PRE_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2A_VITAL of DL2A is
   for VITAL_ACT
   end for;
end CFG_DL2A_VITAL;


----- CELL DL2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2B : entity is TRUE;
end DL2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  H,  x,  x,  S ),
    ( L,  x,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  L,  x,  H ),
    ( U,  x,  x,  x,  H,  H ),
    ( L,  U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Tviol_CLR_G_posedge or Pviol_PRE or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL2B_QN_tab,
        DataIn => (
               CLR_ipd, PRE_ipd, G_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2B_VITAL of DL2B is
   for VITAL_ACT
   end for;
end CFG_DL2B_VITAL;


----- CELL DL2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2C : entity is TRUE;
end DL2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  x,  H ),
    ( H,  H,  x,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  H ),
    ( x,  L,  L,  L,  x,  L ),
    ( U,  x,  x,  x,  L,  L ),
    ( H,  x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Tviol_CLR_G_posedge or Pviol_PRE or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL2C_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2C_VITAL of DL2C is
   for VITAL_ACT
   end for;
end CFG_DL2C_VITAL;


----- CELL DL2D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2D : entity is TRUE;
end DL2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2D_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  x,  L,  x,  S ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  H,  x,  H ),
    ( U,  x,  x,  x,  H,  H ),
    ( L,  U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL2D_QN_tab,
        DataIn => (
               CLR_ipd, PRE_ipd, D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2D_VITAL of DL2D is
   for VITAL_ACT
   end for;
end CFG_DL2D_VITAL;


----- CELL DLC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC : entity is TRUE;
end DLC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC_Q_tab,
        DataIn => (
               CLR_ipd, D_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC_VITAL of DLC is
   for VITAL_ACT
   end for;
end CFG_DLC_VITAL;


----- CELL DLC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1 : entity is TRUE;
end DLC1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1_Q_tab : VitalStateTableType := (
    ( L,  H,  x,  x,  L ),
    ( H,  H,  L,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  L ),
    ( x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1_Q_tab,
        DataIn => (
               D_ipd, G_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1_VITAL of DLC1 is
   for VITAL_ACT
   end for;
end CFG_DLC1_VITAL;


----- CELL DLC1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1A : entity is TRUE;
end DLC1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1A_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  L ),
    ( L,  H,  L,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  L ),
    ( x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1A_Q_tab,
        DataIn => (
               G_ipd, D_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1A_VITAL of DLC1A is
   for VITAL_ACT
   end for;
end CFG_DLC1A_VITAL;


----- CELL DLC1F -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1F is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1F : entity is TRUE;
end DLC1F;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1F is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1F_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( L,  x,  L,  x,  S ),
    ( H,  x,  x,  x,  H ),
    ( x,  L,  H,  x,  H ),
    ( U,  x,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLC1F_QN_tab,
        DataIn => (
               CLR_ipd, D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1F_VITAL of DLC1F is
   for VITAL_ACT
   end for;
end CFG_DLC1F_VITAL;


----- CELL DLC1G -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1G is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1G : entity is TRUE;
end DLC1G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1G is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1G_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H ),
    ( H,  L,  x,  x,  S ),
    ( x,  H,  x,  x,  H ),
    ( x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLC1G_QN_tab,
        DataIn => (
               G_ipd, CLR_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1G_VITAL of DLC1G is
   for VITAL_ACT
   end for;
end CFG_DLC1G_VITAL;


----- CELL DLCA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCA : entity is TRUE;
end DLCA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLCA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLCA_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  L,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLCA_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLCA_VITAL of DLCA is
   for VITAL_ACT
   end for;
end CFG_DLCA_VITAL;


----- CELL DLE -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE : entity is TRUE;
end DLE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( x,  L,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_negedge,
          TimingData              => Tmkr_D_E_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_negedge,
          SetupLow                => tsetup_D_E_noedge_negedge,
          HoldHigh                => thold_D_E_noedge_negedge,
          HoldLow                 => thold_D_E_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_E_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_D_E_negedge or Pviol_E or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE_Q_tab,
        DataIn => (
               D_ipd, G_ipd, E_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE_VITAL of DLE is
   for VITAL_ACT
   end for;
end CFG_DLE_VITAL;


----- CELL DLE1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE1D : entity is TRUE;
end DLE1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE1D_QN_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H ),
    ( L,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLE1D_QN_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (E_ipd'last_event, tpd_E_QN, TRUE),
                 2 => (G_ipd'last_event, tpd_G_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE1D_VITAL of DLE1D is
   for VITAL_ACT
   end for;
end CFG_DLE1D_VITAL;


----- CELL DLE2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE2B : entity is TRUE;
end DLE2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT G_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_E_posedge,
          TimingData              => Tmkr_CLR_E_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_E_posedge_posedge,
          Removal                 => thold_CLR_E_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            =>
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT G_ipd)) /= '0',
          HeaderMsg               => InstancePath &"/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          HeaderMsg               => InstancePath &"/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE2B_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, E_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE2B_VITAL of DLE2B is
   for VITAL_ACT
   end for;
end CFG_DLE2B_VITAL;


----- CELL DLE2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE2C : entity is TRUE;
end DLE2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE2C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR E_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR G_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_E_posedge,
          TimingData              => Tmkr_CLR_E_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_E_negedge_posedge,
          Removal                 => thold_CLR_E_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR G_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR E_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE2C_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE2C_VITAL of DLE2C is
   for VITAL_ACT
   end for;
end CFG_DLE2C_VITAL;


----- CELL DLE3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE3B : entity is TRUE;
end DLE3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE3B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  H ),
    ( x,  x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR E_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR G_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_E_posedge,
          TimingData              => Tmkr_PRE_E_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_E_negedge_posedge,
          Removal                 => thold_PRE_E_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR G_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR E_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_E or Pviol_PRE or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE3B_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE3B_VITAL of DLE3B is
   for VITAL_ACT
   end for;
end CFG_DLE3B_VITAL;


----- CELL DLE3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE3C : entity is TRUE;
end DLE3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE3C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  H,  x,  S ),
    ( x,  H,  x,  H,  x,  S ),
    ( x,  x,  x,  L,  x,  H ),
    ( x,  x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR E_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR G_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_E_posedge,
          TimingData              => Tmkr_PRE_E_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_E_posedge_posedge,
          Removal                 => thold_PRE_E_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR G_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR E_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_E or Pviol_PRE or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE3C_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE3C_VITAL of DLE3C is
   for VITAL_ACT
   end for;
end CFG_DLE3C_VITAL;


----- CELL DLEA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLEA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLEA : entity is TRUE;
end DLEA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLEA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DF1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_E_posedge or Tviol_D_G_negedge or Pviol_E or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               E_ipd, D_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLEA_VITAL of DLEA is
   for VITAL_ACT
   end for;
end CFG_DLEA_VITAL;


----- CELL DLEB -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLEB is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLEB : entity is TRUE;
end DLEB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLEB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_E_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DF1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_negedge,
          TimingData              => Tmkr_D_E_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_negedge,
          SetupLow                => tsetup_D_E_noedge_negedge,
          HoldHigh                => thold_D_E_noedge_negedge,
          HoldLow                 => thold_D_E_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_E_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_E_negedge or Pviol_E or Tviol_D_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               G_ipd, D_ipd, E_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLEB_VITAL of DLEB is
   for VITAL_ACT
   end for;
end CFG_DLEB_VITAL;


----- CELL DLEC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLEC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLEC : entity is TRUE;
end DLEC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLEC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLEC_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLEC_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLEC_VITAL of DLEC is
   for VITAL_ACT
   end for;
end CFG_DLEC_VITAL;


----- CELL DLM -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM : entity is TRUE;
end DLM;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  H,  x,  H ),
    ( x,  L,  L,  H,  x,  L ),
    ( x,  H,  L,  H,  x,  H ),
    ( x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_negedge,
          TimingData              => Tmkr_A_G_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_negedge,
          SetupLow                => tsetup_A_G_noedge_negedge,
          HoldHigh                => thold_A_G_noedge_negedge,
          HoldLow                 => thold_A_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_negedge,
          TimingData              => Tmkr_B_G_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_negedge,
          SetupLow                => tsetup_B_G_noedge_negedge,
          HoldHigh                => thold_B_G_noedge_negedge,
          HoldLow                 => thold_B_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_negedge,
          TimingData              => Tmkr_S_G_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_negedge,
          SetupLow                => tsetup_S_G_noedge_negedge,
          HoldHigh                => thold_S_G_noedge_negedge,
          HoldLow                 => thold_S_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_negedge or Tviol_B_G_negedge or Tviol_S_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM_Q_tab,
        DataIn => (
               B_ipd, A_ipd, S_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM_VITAL of DLM is
   for VITAL_ACT
   end for;
end CFG_DLM_VITAL;


----- CELL DLM2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM2 : entity is TRUE;
end DLM2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM2_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  x,  L ),
    ( x,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_negedge,
          TimingData              => Tmkr_A_G_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_negedge,
          SetupLow                => tsetup_A_G_noedge_negedge,
          HoldHigh                => thold_A_G_noedge_negedge,
          HoldLow                 => thold_A_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_negedge,
          TimingData              => Tmkr_B_G_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_negedge,
          SetupLow                => tsetup_B_G_noedge_negedge,
          HoldHigh                => thold_B_G_noedge_negedge,
          HoldLow                 => thold_B_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_negedge,
          TimingData              => Tmkr_S_G_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_negedge,
          SetupLow                => tsetup_S_G_noedge_negedge,
          HoldHigh                => thold_S_G_noedge_negedge,
          HoldLow                 => thold_S_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_negedge or Tviol_B_G_negedge or Tviol_S_G_negedge or Pviol_CLR or Tviol_CLR_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM2_Q_tab,
        DataIn => (
               CLR_ipd, B_ipd, A_ipd, S_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 4 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM2_VITAL of DLM2 is
   for VITAL_ACT
   end for;
end CFG_DLM2_VITAL;


----- CELL DLM2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM2B : entity is TRUE;
end DLM2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_posedge,
          TimingData              => Tmkr_A_G_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_posedge,
          SetupLow                => tsetup_A_G_noedge_posedge,
          HoldHigh                => thold_A_G_noedge_posedge,
          HoldLow                 => thold_A_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_posedge,
          TimingData              => Tmkr_B_G_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_posedge,
          SetupLow                => tsetup_B_G_noedge_posedge,
          HoldHigh                => thold_B_G_noedge_posedge,
          HoldLow                 => thold_B_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_posedge,
          TimingData              => Tmkr_S_G_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_posedge,
          SetupLow                => tsetup_S_G_noedge_posedge,
          HoldHigh                => thold_S_G_noedge_posedge,
          HoldLow                 => thold_S_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_posedge or Tviol_B_G_posedge or Tviol_CLR_G_posedge or Tviol_S_G_posedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM2B_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, B_ipd, A_ipd, S_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 4 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM2B_VITAL of DLM2B is
   for VITAL_ACT
   end for;
end CFG_DLM2B_VITAL;


----- CELL DLM3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM3 : entity is TRUE;
end DLM3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_negedge,
          TimingData              => Tmkr_D0_G_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_negedge,
          SetupLow                => tsetup_D0_G_noedge_negedge,
          HoldHigh                => thold_D0_G_noedge_negedge,
          HoldLow                 => thold_D0_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_negedge,
          TimingData              => Tmkr_D1_G_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_negedge,
          SetupLow                => tsetup_D1_G_noedge_negedge,
          HoldHigh                => thold_D1_G_noedge_negedge,
          HoldLow                 => thold_D1_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_negedge,
          TimingData              => Tmkr_D2_G_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_negedge,
          SetupLow                => tsetup_D2_G_noedge_negedge,
          HoldHigh                => thold_D2_G_noedge_negedge,
          HoldLow                 => thold_D2_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_negedge,
          TimingData              => Tmkr_D3_G_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_negedge,
          SetupLow                => tsetup_D3_G_noedge_negedge,
          HoldHigh                => thold_D3_G_noedge_negedge,
          HoldLow                 => thold_D3_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_negedge,
          TimingData              => Tmkr_S0_G_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_negedge,
          SetupLow                => tsetup_S0_G_noedge_negedge,
          HoldHigh                => thold_S0_G_noedge_negedge,
          HoldLow                 => thold_S0_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_G_negedge,
          TimingData              => Tmkr_S1_G_negedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_G_noedge_negedge,
          SetupLow                => tsetup_S1_G_noedge_negedge,
          HoldHigh                => thold_S1_G_noedge_negedge,
          HoldLow                 => thold_S1_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_negedge or Tviol_D2_G_negedge or Tviol_D3_G_negedge or Tviol_S0_G_negedge or Tviol_S1_G_negedge or Tviol_D1_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM3_Q_tab,
        DataIn => (
               D3_ipd, D2_ipd, D1_ipd, D0_ipd, S1_ipd, S0_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 6 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM3_VITAL of DLM3 is
   for VITAL_ACT
   end for;
end CFG_DLM3_VITAL;


----- CELL DLM3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM3A : entity is TRUE;
end DLM3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM3A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_posedge,
          TimingData              => Tmkr_D0_G_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_posedge,
          SetupLow                => tsetup_D0_G_noedge_posedge,
          HoldHigh                => thold_D0_G_noedge_posedge,
          HoldLow                 => thold_D0_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_posedge,
          TimingData              => Tmkr_D1_G_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_posedge,
          SetupLow                => tsetup_D1_G_noedge_posedge,
          HoldHigh                => thold_D1_G_noedge_posedge,
          HoldLow                 => thold_D1_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_posedge,
          TimingData              => Tmkr_D2_G_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_posedge,
          SetupLow                => tsetup_D2_G_noedge_posedge,
          HoldHigh                => thold_D2_G_noedge_posedge,
          HoldLow                 => thold_D2_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_posedge,
          TimingData              => Tmkr_D3_G_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_posedge,
          SetupLow                => tsetup_D3_G_noedge_posedge,
          HoldHigh                => thold_D3_G_noedge_posedge,
          HoldLow                 => thold_D3_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_posedge,
          TimingData              => Tmkr_S0_G_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_posedge,
          SetupLow                => tsetup_S0_G_noedge_posedge,
          HoldHigh                => thold_S0_G_noedge_posedge,
          HoldLow                 => thold_S0_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_G_posedge,
          TimingData              => Tmkr_S1_G_posedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_G_noedge_posedge,
          SetupLow                => tsetup_S1_G_noedge_posedge,
          HoldHigh                => thold_S1_G_noedge_posedge,
          HoldLow                 => thold_S1_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_posedge or Tviol_S0_G_posedge or Tviol_S1_G_posedge or Tviol_D1_G_posedge or Tviol_D2_G_posedge or Tviol_D3_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM3A_Q_tab,
        DataIn => (
               G_ipd, D3_ipd, D2_ipd, D1_ipd, D0_ipd, S1_ipd, S0_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 6 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM3A_VITAL of DLM3A is
   for VITAL_ACT
   end for;
end CFG_DLM3A_VITAL;


----- CELL DLM4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM4 : entity is TRUE;
end DLM4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM4_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_negedge,
          TimingData              => Tmkr_D0_G_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_negedge,
          SetupLow                => tsetup_D0_G_noedge_negedge,
          HoldHigh                => thold_D0_G_noedge_negedge,
          HoldLow                 => thold_D0_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_negedge,
          TimingData              => Tmkr_D1_G_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_negedge,
          SetupLow                => tsetup_D1_G_noedge_negedge,
          HoldHigh                => thold_D1_G_noedge_negedge,
          HoldLow                 => thold_D1_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_negedge,
          TimingData              => Tmkr_D2_G_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_negedge,
          SetupLow                => tsetup_D2_G_noedge_negedge,
          HoldHigh                => thold_D2_G_noedge_negedge,
          HoldLow                 => thold_D2_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_negedge,
          TimingData              => Tmkr_D3_G_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_negedge,
          SetupLow                => tsetup_D3_G_noedge_negedge,
          HoldHigh                => thold_D3_G_noedge_negedge,
          HoldLow                 => thold_D3_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_negedge,
          TimingData              => Tmkr_S0_G_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_negedge,
          SetupLow                => tsetup_S0_G_noedge_negedge,
          HoldHigh                => thold_S0_G_noedge_negedge,
          HoldLow                 => thold_S0_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_G_negedge,
          TimingData              => Tmkr_S10_G_negedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_G_noedge_negedge,
          SetupLow                => tsetup_S10_G_noedge_negedge,
          HoldHigh                => thold_S10_G_noedge_negedge,
          HoldLow                 => thold_S10_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_G_negedge,
          TimingData              => Tmkr_S11_G_negedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_G_noedge_negedge,
          SetupLow                => tsetup_S11_G_noedge_negedge,
          HoldHigh                => thold_S11_G_noedge_negedge,
          HoldLow                 => thold_S11_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_negedge or Tviol_D2_G_negedge or Tviol_D3_G_negedge or Tviol_S0_G_negedge or Tviol_D1_G_negedge or Tviol_S10_G_negedge or Pviol_G or Tviol_S11_G_negedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM4_Q_tab,
        DataIn => (
               D3_ipd, D2_ipd, D1_ipd, D0_ipd, S11_ipd, S10_ipd, S0_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S10_ipd'last_event, tpd_S10_Q, TRUE),
                 6 => (S11_ipd'last_event, tpd_S11_Q, TRUE),
                 7 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM4_VITAL of DLM4 is
   for VITAL_ACT
   end for;
end CFG_DLM4_VITAL;


----- CELL DLM4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM4A : entity is TRUE;
end DLM4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM4A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_posedge,
          TimingData              => Tmkr_D0_G_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_posedge,
          SetupLow                => tsetup_D0_G_noedge_posedge,
          HoldHigh                => thold_D0_G_noedge_posedge,
          HoldLow                 => thold_D0_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_posedge,
          TimingData              => Tmkr_D1_G_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_posedge,
          SetupLow                => tsetup_D1_G_noedge_posedge,
          HoldHigh                => thold_D1_G_noedge_posedge,
          HoldLow                 => thold_D1_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_posedge,
          TimingData              => Tmkr_D2_G_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_posedge,
          SetupLow                => tsetup_D2_G_noedge_posedge,
          HoldHigh                => thold_D2_G_noedge_posedge,
          HoldLow                 => thold_D2_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_posedge,
          TimingData              => Tmkr_D3_G_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_posedge,
          SetupLow                => tsetup_D3_G_noedge_posedge,
          HoldHigh                => thold_D3_G_noedge_posedge,
          HoldLow                 => thold_D3_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_posedge,
          TimingData              => Tmkr_S0_G_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_posedge,
          SetupLow                => tsetup_S0_G_noedge_posedge,
          HoldHigh                => thold_S0_G_noedge_posedge,
          HoldLow                 => thold_S0_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_G_posedge,
          TimingData              => Tmkr_S10_G_posedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_G_noedge_posedge,
          SetupLow                => tsetup_S10_G_noedge_posedge,
          HoldHigh                => thold_S10_G_noedge_posedge,
          HoldLow                 => thold_S10_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_G_posedge,
          TimingData              => Tmkr_S11_G_posedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_G_noedge_posedge,
          SetupLow                => tsetup_S11_G_noedge_posedge,
          HoldHigh                => thold_S11_G_noedge_posedge,
          HoldLow                 => thold_S11_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_posedge or Tviol_S0_G_posedge or Tviol_D1_G_posedge or Tviol_D2_G_posedge or Tviol_D3_G_posedge or Tviol_S10_G_posedge or Tviol_S11_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM4A_Q_tab,
        DataIn => (
               G_ipd, D3_ipd, D2_ipd, D1_ipd, D0_ipd, S11_ipd, S10_ipd, S0_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S10_ipd'last_event, tpd_S10_Q, TRUE),
                 6 => (S11_ipd'last_event, tpd_S11_Q, TRUE),
                 7 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM4A_VITAL of DLM4A is
   for VITAL_ACT
   end for;
end CFG_DLM4A_VITAL;


----- CELL DLM8A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM8A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S00_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S01_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S00_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S00_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S01_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S01_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S00                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S01                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM8A : entity is TRUE;
end DLM8A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM8A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S00_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S01_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S00_ipd, S00, tipd_S00);
   VitalWireDelay (S01_ipd, S01, tipd_S01);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S00_ipd, S01_ipd, S10_ipd, S11_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S00_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S00_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S01_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S01_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 9);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM8A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  H,  H,  H,  H,  x,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  H,  x,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  H,  x,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  x,  x,  x,  L,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  x,  x,  x,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  L,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  x,  H,  x,  H,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  H,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  x,  H,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  H,  H,  L,  L,  x,  x,  H,  x,  H ),
    ( H,  x,  x,  H,  x,  L,  L,  L,  x,  H,  x,  H ),
    ( H,  x,  x,  H,  x,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  L,  L,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  H,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  x,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  x,  H,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  x,  L,  x,  x,  H,  x,  H,  H,  H,  x,  L ),
    ( x,  x,  L,  x,  x,  x,  H,  H,  H,  H,  x,  L ),
    ( x,  x,  x,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  x,  x,  x,  L,  L,  L,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_negedge,
          TimingData              => Tmkr_D0_G_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_negedge,
          SetupLow                => tsetup_D0_G_noedge_negedge,
          HoldHigh                => thold_D0_G_noedge_negedge,
          HoldLow                 => thold_D0_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_negedge,
          TimingData              => Tmkr_D1_G_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_negedge,
          SetupLow                => tsetup_D1_G_noedge_negedge,
          HoldHigh                => thold_D1_G_noedge_negedge,
          HoldLow                 => thold_D1_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd ))
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_negedge,
          TimingData              => Tmkr_D2_G_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_negedge,
          SetupLow                => tsetup_D2_G_noedge_negedge,
          HoldHigh                => thold_D2_G_noedge_negedge,
          HoldLow                 => thold_D2_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_negedge,
          TimingData              => Tmkr_D3_G_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_negedge,
          SetupLow                => tsetup_D3_G_noedge_negedge,
          HoldHigh                => thold_D3_G_noedge_negedge,
          HoldLow                 => thold_D3_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd ))
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S00_G_negedge,
          TimingData              => Tmkr_S00_G_negedge,
          TestSignal              => S00_ipd,
          TestSignalName          => "S00",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S00_G_noedge_negedge,
          SetupLow                => tsetup_S00_G_noedge_negedge,
          HoldHigh                => thold_S00_G_noedge_negedge,
          HoldLow                 => thold_S00_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S01_G_negedge,
          TimingData              => Tmkr_S01_G_negedge,
          TestSignal              => S01_ipd,
          TestSignalName          => "S01",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S01_G_noedge_negedge,
          SetupLow                => tsetup_S01_G_noedge_negedge,
          HoldHigh                => thold_S01_G_noedge_negedge,
          HoldLow                 => thold_S01_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_G_negedge,
          TimingData              => Tmkr_S10_G_negedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_G_noedge_negedge,
          SetupLow                => tsetup_S10_G_noedge_negedge,
          HoldHigh                => thold_S10_G_noedge_negedge,
          HoldLow                 => thold_S10_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_G_negedge,
          TimingData              => Tmkr_S11_G_negedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_G_noedge_negedge,
          SetupLow                => tsetup_S11_G_noedge_negedge,
          HoldHigh                => thold_S11_G_noedge_negedge,
          HoldLow                 => thold_S11_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM8A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_negedge or Tviol_D2_G_negedge or Tviol_D3_G_negedge or Tviol_S00_G_negedge or Tviol_S01_G_negedge or Pviol_CLR or Tviol_D1_G_negedge or Tviol_S10_G_negedge or Tviol_CLR_G_negedge or Pviol_G or Tviol_S11_G_negedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM8A_Q_tab,
        DataIn => (
               CLR_ipd, D2_ipd, D3_ipd, D0_ipd, D1_ipd, S11_ipd, S10_ipd, S01_ipd, S00_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S00_ipd'last_event, tpd_S00_Q, TRUE),
                 5 => (S01_ipd'last_event, tpd_S01_Q, TRUE),
                 6 => (S10_ipd'last_event, tpd_S10_Q, TRUE),
                 7 => (S11_ipd'last_event, tpd_S11_Q, TRUE),
                 8 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 9 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM8A_VITAL of DLM8A is
   for VITAL_ACT
   end for;
end CFG_DLM8A_VITAL;


----- CELL DLM8B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM8B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S00_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S01_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S00_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S00_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S01_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S01_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S00                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S01                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM8B : entity is TRUE;
end DLM8B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of DLM8B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S00_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S01_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S00_ipd, S00, tipd_S00);
   VitalWireDelay (S01_ipd, S01, tipd_S01);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S00_ipd, S01_ipd, S10_ipd, S11_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S00_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S00_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S01_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S01_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 9);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM8B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  x,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  x,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  L,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  x,  L,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  L,  x,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  x,  L,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  L,  x,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  x,  L,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  x,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  L,  x,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  x,  L,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  x,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  x,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  x,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  x,  L,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  x,  L,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  x,  L,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  x,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  L,  x,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  x,  L,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_posedge,
          TimingData              => Tmkr_D0_G_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_posedge,
          SetupLow                => tsetup_D0_G_noedge_posedge,
          HoldHigh                => thold_D0_G_noedge_posedge,
          HoldLow                 => thold_D0_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_posedge,
          TimingData              => Tmkr_D1_G_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_posedge,
          SetupLow                => tsetup_D1_G_noedge_posedge,
          HoldHigh                => thold_D1_G_noedge_posedge,
          HoldLow                 => thold_D1_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd ))
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_posedge,
          TimingData              => Tmkr_D2_G_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_posedge,
          SetupLow                => tsetup_D2_G_noedge_posedge,
          HoldHigh                => thold_D2_G_noedge_posedge,
          HoldLow                 => thold_D2_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S00_ipd AND S01_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_posedge,
          TimingData              => Tmkr_D3_G_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_posedge,
          SetupLow                => tsetup_D3_G_noedge_posedge,
          HoldHigh                => thold_D3_G_noedge_posedge,
          HoldLow                 => thold_D3_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT ( S00_ipd AND S01_ipd ))
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S00_G_posedge,
          TimingData              => Tmkr_S00_G_posedge,
          TestSignal              => S00_ipd,
          TestSignalName          => "S00",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S00_G_noedge_posedge,
          SetupLow                => tsetup_S00_G_noedge_posedge,
          HoldHigh                => thold_S00_G_noedge_posedge,
          HoldLow                 => thold_S00_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S01_G_posedge,
          TimingData              => Tmkr_S01_G_posedge,
          TestSignal              => S01_ipd,
          TestSignalName          => "S01",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S01_G_noedge_posedge,
          SetupLow                => tsetup_S01_G_noedge_posedge,
          HoldHigh                => thold_S01_G_noedge_posedge,
          HoldLow                 => thold_S01_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_G_posedge,
          TimingData              => Tmkr_S10_G_posedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_G_noedge_posedge,
          SetupLow                => tsetup_S10_G_noedge_posedge,
          HoldHigh                => thold_S10_G_noedge_posedge,
          HoldLow                 => thold_S10_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_G_posedge,
          TimingData              => Tmkr_S11_G_posedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_G_noedge_posedge,
          SetupLow                => tsetup_S11_G_noedge_posedge,
          HoldHigh                => thold_S11_G_noedge_posedge,
          HoldLow                 => thold_S11_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM8B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_posedge or Tviol_D1_G_posedge or Tviol_D2_G_posedge or Tviol_D3_G_posedge or Tviol_S10_G_posedge or Tviol_CLR_G_posedge or Tviol_S11_G_posedge or Tviol_S00_G_posedge or Pviol_G or Pviol_CLR or Tviol_S01_G_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM8B_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, D2_ipd, D3_ipd, D0_ipd, D1_ipd, S11_ipd, S10_ipd, S01_ipd, S00_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S00_ipd'last_event, tpd_S00_Q, TRUE),
                 5 => (S01_ipd'last_event, tpd_S01_Q, TRUE),
                 6 => (S10_ipd'last_event, tpd_S10_Q, TRUE),
                 7 => (S11_ipd'last_event, tpd_S11_Q, TRUE),
                 8 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 9 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM8B_VITAL of DLM8B is
   for VITAL_ACT
   end for;
end CFG_DLM8B_VITAL;


----- CELL DLMA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLMA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLMA : entity is TRUE;
end DLMA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLMA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLMA_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  x,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L ),
    ( L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_posedge,
          TimingData              => Tmkr_A_G_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_posedge,
          SetupLow                => tsetup_A_G_noedge_posedge,
          HoldHigh                => thold_A_G_noedge_posedge,
          HoldLow                 => thold_A_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_posedge,
          TimingData              => Tmkr_B_G_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_posedge,
          SetupLow                => tsetup_B_G_noedge_posedge,
          HoldHigh                => thold_B_G_noedge_posedge,
          HoldLow                 => thold_B_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_posedge,
          TimingData              => Tmkr_S_G_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_posedge,
          SetupLow                => tsetup_S_G_noedge_posedge,
          HoldHigh                => thold_S_G_noedge_posedge,
          HoldLow                 => thold_S_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_posedge or Tviol_B_G_posedge or Tviol_S_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLMA_Q_tab,
        DataIn => (
               G_ipd, B_ipd, A_ipd, S_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLMA_VITAL of DLMA is
   for VITAL_ACT
   end for;
end CFG_DLMA_VITAL;


----- CELL DLME1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLME1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_A_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_A_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_B_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_B_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_S_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLME1A : entity is TRUE;
end DLME1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLME1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_A_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  H,  H,  x,  x,  H ),
    ( L,  L,  H,  x,  H,  x,  H ),
    ( L,  L,  x,  L,  L,  x,  L ),
    ( L,  L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_posedge,
          TimingData              => Tmkr_A_G_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_posedge,
          SetupLow                => tsetup_A_G_noedge_posedge,
          HoldHigh                => thold_A_G_noedge_posedge,
          HoldLow                 => thold_A_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_A_E_posedge,
          TimingData              => Tmkr_A_E_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_E_noedge_posedge,
          SetupLow                => tsetup_A_E_noedge_posedge,
          HoldHigh                => thold_A_E_noedge_posedge,
          HoldLow                 => thold_A_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_posedge,
          TimingData              => Tmkr_B_G_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_posedge,
          SetupLow                => tsetup_B_G_noedge_posedge,
          HoldHigh                => thold_B_G_noedge_posedge,
          HoldLow                 => thold_B_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR (NOT S_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_E_posedge,
          TimingData              => Tmkr_B_E_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_E_noedge_posedge,
          SetupLow                => tsetup_B_E_noedge_posedge,
          HoldHigh                => thold_B_E_noedge_posedge,
          HoldLow                 => thold_B_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_posedge,
          TimingData              => Tmkr_S_G_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_posedge,
          SetupLow                => tsetup_S_G_noedge_posedge,
          HoldHigh                => thold_S_G_noedge_posedge,
          HoldLow                 => thold_S_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_E_posedge,
          TimingData              => Tmkr_S_E_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_E_noedge_posedge,
          SetupLow                => tsetup_S_E_noedge_posedge,
          HoldHigh                => thold_S_E_noedge_posedge,
          HoldLow                 => thold_S_E_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_posedge or Pviol_E or Tviol_A_E_posedge or Tviol_B_G_posedge or Tviol_B_E_posedge or Tviol_S_G_posedge or Tviol_S_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLME1A_Q_tab,
        DataIn => (
               G_ipd, E_ipd, B_ipd, A_ipd, S_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 4 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLME1A_VITAL of DLME1A is
   for VITAL_ACT
   end for;
end CFG_DLME1A_VITAL;


----- CELL DLP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1 : entity is TRUE;
end DLP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  H,  x,  x,  H ),
    ( x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1_Q_tab,
        DataIn => (
               D_ipd, PRE_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1_VITAL of DLP1 is
   for VITAL_ACT
   end for;
end CFG_DLP1_VITAL;


----- CELL DLP1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1A : entity is TRUE;
end DLP1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  H ),
    ( x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1A_Q_tab,
        DataIn => (
               G_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1A_VITAL of DLP1A is
   for VITAL_ACT
   end for;
end CFG_DLP1A_VITAL;


----- CELL DLP1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1B : entity is TRUE;
end DLP1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1B_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  x,  x,  H ),
    ( x,  H,  L,  x,  S ),
    ( x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1B_Q_tab,
        DataIn => (
               D_ipd, PRE_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1B_VITAL of DLP1B is
   for VITAL_ACT
   end for;
end CFG_DLP1B_VITAL;


----- CELL DLP1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1C : entity is TRUE;
end DLP1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1C_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  H,  x,  S ),
    ( x,  x,  L,  x,  H ),
    ( x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1C_Q_tab,
        DataIn => (
               G_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1C_VITAL of DLP1C is
   for VITAL_ACT
   end for;
end CFG_DLP1C_VITAL;


----- CELL DLP1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1D : entity is TRUE;
end DLP1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1D_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  H,  H,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLP1D_QN_tab,
        DataIn => (
               PRE_ipd, D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1D_VITAL of DLP1D is
   for VITAL_ACT
   end for;
end CFG_DLP1D_VITAL;


----- CELL DLP1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1E : entity is TRUE;
end DLP1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLP1E_QN_tab,
        DataIn => (
               PRE_ipd, G_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1E_VITAL of DLP1E is
   for VITAL_ACT
   end for;
end CFG_DLP1E_VITAL;


----- CELL FA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity FA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of FA1A : entity is TRUE;
end FA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of FA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS S_zd : STD_LOGIC is Results(1);
   ALIAS CO_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE S_GlitchData	: VitalGlitchDataType;
   VARIABLE CO_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      S_zd :=
       (((NOT A_ipd)) AND ((((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND
         (CI_ipd) AND ((NOT A_ipd))) OR ((CI_ipd) AND (B_ipd) AND (A_ipd)))
         AND (CI_ipd)) OR (((NOT A_ipd)) AND (B_ipd) AND ((NOT CI_ipd))) OR
         ((A_ipd) AND ((((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND
         (CI_ipd) AND ((NOT A_ipd))) OR ((CI_ipd) AND (B_ipd) AND (A_ipd)))
         AND ((NOT CI_ipd))) OR ((A_ipd) AND (B_ipd) AND (CI_ipd));
      CO_zd :=
       (((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND (CI_ipd)) OR 
       ((CI_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_FA1A_VITAL of FA1A is
   for VITAL_ACT
   end for;
end CFG_FA1A_VITAL;


----- CELL FA1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity FA1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of FA1B : entity is TRUE;
end FA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of FA1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS S_zd : STD_LOGIC is Results(1);
   ALIAS CO_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE S_GlitchData	: VitalGlitchDataType;
   VARIABLE CO_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      S_zd :=
       ((((((CI_ipd) AND ((NOT B_ipd)) AND (A_ipd)) OR ((((CI_ipd) AND
         (B_ipd)) OR ((NOT B_ipd))) AND ((NOT A_ipd)))) AND (CI_ipd)) OR
         ((B_ipd) AND ((NOT CI_ipd)))) AND (A_ipd)) OR ((((B_ipd) AND
         (CI_ipd)) OR ((((CI_ipd) AND ((NOT B_ipd)) AND (A_ipd)) OR
         ((((CI_ipd) AND (B_ipd)) OR ((NOT B_ipd))) AND ((NOT A_ipd)))) AND
         ((NOT CI_ipd)))) AND ((NOT A_ipd)));
      CO_zd :=
       ((CI_ipd) AND ((NOT B_ipd))) OR ((CI_ipd) AND ((NOT A_ipd)))
         OR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_FA1B_VITAL of FA1B is
   for VITAL_ACT
   end for;
end CFG_FA1B_VITAL;


----- CELL FA2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity FA2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of FA2A : entity is TRUE;
end FA2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of FA2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS S_zd : STD_LOGIC is Results(1);
   ALIAS CO_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE S_GlitchData	: VitalGlitchDataType;
   VARIABLE CO_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      S_zd :=
       (((NOT ((A1_ipd) OR (A0_ipd)))) AND ((((A1_ipd) OR (A0_ipd)) AND
         ((NOT B_ipd))) OR (((NOT B_ipd)) AND (CI_ipd) AND ((NOT ((A1_ipd) OR
         (A0_ipd))))) OR ((CI_ipd) AND (B_ipd) AND ((A1_ipd) OR (A0_ipd))))
         AND (CI_ipd)) OR (((NOT ((A1_ipd) OR (A0_ipd)))) AND (B_ipd) AND
         ((NOT CI_ipd))) OR (((A1_ipd) OR (A0_ipd)) AND ((((A1_ipd) OR
         (A0_ipd)) AND ((NOT B_ipd))) OR (((NOT B_ipd)) AND (CI_ipd) AND
         ((NOT ((A1_ipd) OR (A0_ipd))))) OR ((CI_ipd) AND (B_ipd) AND
         ((A1_ipd) OR (A0_ipd)))) AND ((NOT CI_ipd))) OR (((A1_ipd) OR
         (A0_ipd)) AND (B_ipd) AND (CI_ipd));
      --CO_zd :=
      -- (((A1_ipd) OR (A0_ipd)) AND ((NOT B_ipd))) OR (((NOT B_ipd)) AND
      --   (CI_ipd) AND ((NOT ((A1_ipd) OR (A0_ipd))))) OR ((CI_ipd) AND
      --   (B_ipd) AND ((A1_ipd) OR (A0_ipd)));
      CO_zd := 
        (((A1_ipd) AND (NOT B_ipd)) OR ((A0_ipd) AND (NOT B_ipd)) OR
         ((A0_ipd) AND (CI_ipd)) OR ((A1_ipd) AND (CI_ipd)) OR
         ((NOT B_ipd) AND (CI_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_S, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_CO, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_FA2A_VITAL of FA2A is
   for VITAL_ACT
   end for;
end CFG_FA2A_VITAL;


----- CELL FECTH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FECTH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
                tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);        -- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FECTH : ENTITY IS TRUE;
	--
end FECTH;

ARCHITECTURE VITAL_ACT OF FECTH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FECTH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FECTH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FECTH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FECTH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FECTH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FECTH_TAB Declaration
		CONSTANT  FECTH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FECTH_TAB
		VitalStateTable (
				StateTable         => FECTH_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FECTH_TAB_Result,
				PreviousDataIn     => PrevData_FECTH_TAB
		);	--End VitalStateTable
		FECTH_TABStateReg(0)     := FECTH_TAB_Result(2);
		LSB(0)                    := FECTH_TAB_Result(1);
		Y_zd                      := LSB(0);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FECTH_VITAL of FECTH is
   for VITAL_ACT
   end for;
end CFG_FECTH_VITAL;
----- CELL FECTL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FECTL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
                tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);        -- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FECTL : ENTITY IS TRUE;
	--
end FECTL;

ARCHITECTURE VITAL_ACT OF FECTL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FECTL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FECTL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FECTL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FECTL_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FECTL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FECTL_TAB Declaration
		CONSTANT  FECTL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FECTL_TAB
		VitalStateTable (
				StateTable         => FECTL_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FECTL_TAB_Result,
				PreviousDataIn     => PrevData_FECTL_TAB
		);	--End VitalStateTable
		FECTL_TABStateReg(0)     := FECTL_TAB_Result(2);
		LSB(0)                    := FECTL_TAB_Result(1);
		Y_zd                      := LSB(0);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FECTL_VITAL of FECTL is
   for VITAL_ACT
   end for;
end CFG_FECTL_VITAL;
----- CELL FECTMH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FECTMH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FECTMH : ENTITY IS TRUE;
	--
end FECTMH;

ARCHITECTURE VITAL_ACT OF FECTMH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    M_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => M_ipd,
				InSig              => M,
				twire              => tipd_M
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, M_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FECTMH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FECTMH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FECTMH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FECTMH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FECTMH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FECTMH_TAB Declaration
		CONSTANT  FECTMH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FECTMH_TAB
		VitalStateTable (
				StateTable         => FECTMH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FECTMH_TAB_Result,
				PreviousDataIn     => PrevData_FECTMH_TAB
		);	--End VitalStateTable
		FECTMH_TABStateReg(0)     := FECTMH_TAB_Result(2);
		LSB(0)                    := FECTMH_TAB_Result(1);
		Y_zd                      := VitalMux2(data1 => PAD_ipd, data0 => LSB(0), dselect => M_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => M_ipd'LAST_EVENT,
							PathDelay       => tpd_M_Y,
							PathCondition   => TRUE
				                      ),
				                 3 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FECTMH_VITAL of FECTMH is
   for VITAL_ACT
   end for;
end CFG_FECTMH_VITAL;
----- CELL FECTML -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FECTML IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FECTML : ENTITY IS TRUE;
	--
end FECTML;

ARCHITECTURE VITAL_ACT OF FECTML IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    M_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => M_ipd,
				InSig              => M,
				twire              => tipd_M
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, M_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FECTML_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FECTML_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FECTML_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FECTML_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FECTML_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FECTML_TAB Declaration
		CONSTANT  FECTML_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
		( '0', '0', '-', '-', '-',  '-',  '0',  '0' ),
		( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
		( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
		( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
		( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '0', '-',  '0',  '0',  '0' ),
		( '0', '-', '-', '-', '1',  '0',  '0',  '0' ),
		( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
		( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
		( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
		( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
		( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FECTML_TAB
		VitalStateTable (
				StateTable         => FECTML_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FECTML_TAB_Result,
				PreviousDataIn     => PrevData_FECTML_TAB
		);	--End VitalStateTable
		FECTML_TABStateReg(0)     := FECTML_TAB_Result(2);
		LSB(0)                    := FECTML_TAB_Result(1);
		Y_zd                      := VitalMux2(data1 => PAD_ipd, data0 => LSB(0), dselect => M_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => M_ipd'LAST_EVENT,
							PathDelay       => tpd_M_Y,
							PathCondition   => TRUE
				                      ),
				                 3 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FECTML_VITAL of FECTML is
   for VITAL_ACT
   end for;
end CFG_FECTML_VITAL;
----- CELL FEPTH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FEPTH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FEPTH : ENTITY IS TRUE;
	--
end FEPTH;

ARCHITECTURE VITAL_ACT OF FEPTH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd 
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FEPTH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FEPTH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FEPTH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FEPTH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FEPTH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FEPTH_TAB Declaration
		CONSTANT  FEPTH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
                ( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
                ( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
                ( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
                ( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
                ( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
                ( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
                ( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FEPTH_TAB
		VitalStateTable (
				StateTable         => FEPTH_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FEPTH_TAB_Result,
				PreviousDataIn     => PrevData_FEPTH_TAB
		);	--End VitalStateTable
		FEPTH_TABStateReg(0)      := FEPTH_TAB_Result(2);
		LSB(0)                    := FEPTH_TAB_Result(1);
		Y_zd                      := LSB(0);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FEPTH_VITAL of FEPTH is
   for VITAL_ACT
   end for;
end CFG_FEPTH_VITAL;
----- CELL FEPTL -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FEPTL IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : OUT     STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FEPTL : ENTITY IS TRUE;
	--
end FEPTL;

ARCHITECTURE VITAL_ACT OF FEPTL IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd 
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FEPTL_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FEPTL_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FEPTL_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FEPTL_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FEPTL_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FEPTL_TAB Declaration
		CONSTANT  FEPTL_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
                ( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
                ( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
                ( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
                ( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
                ( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
                ( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
                ( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FEPTL_TAB
		VitalStateTable (
				StateTable         => FEPTL_TAB,
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FEPTL_TAB_Result,
				PreviousDataIn     => PrevData_FEPTL_TAB
		);	--End VitalStateTable
		FEPTL_TABStateReg(0)      := FEPTL_TAB_Result(2);
		LSB(0)                    := FEPTL_TAB_Result(1);
		Y_zd                      := LSB(0);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FEPTL_VITAL of FEPTL is
   for VITAL_ACT
   end for;
end CFG_FEPTL_VITAL;
----- CELL FEPTMH -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FEPTMH IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FEPTMH : ENTITY IS TRUE;
	--
end FEPTMH;

ARCHITECTURE VITAL_ACT OF FEPTMH IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    M_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => M_ipd,
				InSig              => M,
				twire              => tipd_M
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, M_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FEPTMH_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FEPTMH_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FEPTMH_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FEPTMH_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FEPTMH_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FEPTMH_TAB Declaration
		CONSTANT  FEPTMH_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
                ( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
                ( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
                ( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
                ( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
                ( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
                ( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
                ( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FEPTMH_TAB
		VitalStateTable (
				StateTable         => FEPTMH_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FEPTMH_TAB_Result,
				PreviousDataIn     => PrevData_FEPTMH_TAB
		);	--End VitalStateTable
		FEPTMH_TABStateReg(0)     := FEPTMH_TAB_Result(2);
		LSB(0)                    := FEPTMH_TAB_Result(1);
		Y_zd                      := VitalMux2(data1 => PAD_ipd, data0 => LSB(0), dselect => M_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => M_ipd'LAST_EVENT,
							PathDelay       => tpd_M_Y,
							PathCondition   => TRUE
				                      ),
				                 3 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FEPTMH_VITAL of FEPTMH is
   for VITAL_ACT
   end for;
end CFG_FEPTMH_VITAL;
----- CELL FEPTML -----
LIBRARY   IEEE;
USE       IEEE.std_logic_1164.all;
USE       IEEE.VITAL_Timing.all;
USE       IEEE.VITAL_Primitives.all;
	
entity FEPTML IS
	GENERIC (
		--
		-- PinToPinDelay Generics Declaration(s)
		tpd_PAD_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input PAD to output Y
		tpd_M_Y              : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input M to output Y
		tpd_IOPCL_PAD        : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output PAD
		tpd_IOPCL_Y          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input IOPCL to output Y
		tpd_CLK_PAD          : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output PAD
		tpd_CLK_Y            : VitalDelayType01 := (1.000 ns, 1.000 ns);	-- Path delay from input CLK to output Y
		tpd_E_PAD            : VitalDelayType01z := (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns); -- Path delay from input E to output PAD

		--
		-- Interconnect Path Delay Generics Declaration(s)
		tipd_CLK             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port CLK
		tipd_D               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port D
		tipd_E               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port E
		tipd_M               : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port M
		tipd_IOPCL           : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port IOPCL
		tipd_ODE             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port ODE
		tipd_PAD             : VitalDelayType01 := (0.000 ns, 0.000 ns);	-- Input wire delay on port PAD
		--
		-- Setup Generics Declaration(s)
		tsetup_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between D and CLK
		tsetup_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Setup Hi time between ODE and CLK
		--
		-- Hold Generics Declaration(s)
		thold_D_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between D and CLK
		thold_ODE_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between ODE and CLK
		thold_IOPCL_CLK_noedge_posedge : VitalDelayType   := 0.000 ns;	-- Hold Hi time between IOPCL and CLK
		--
		-- Recovery Generics Declaration(s)
		trecovery_IOPCL_CLK_posedge_posedge : VitalDelayType   := 0.000 ns;	-- Recovery time between IOPCL and CLK
		--
		-- Period Check Generics Declaration(s)
		tperiod_CLK_posedge          : VitalDelayType   := 0.000 ns;	-- Minimum period time for CLK
		tpw_CLK_posedge      : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for CLK
		tpw_CLK_negedge      : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for CLK
		tperiod_IOPCL        : VitalDelayType   := 0.000 ns;	-- Minimum period time for IOPCL
		tpw_IOPCL_posedge    : VitalDelayType   := 0.000 ns;	-- Minimum high pulse width for IOPCL
		tpw_IOPCL_negedge    : VitalDelayType   := 0.000 ns;	-- Minimum low pulse width for IOPCL
		--
		-- InstancePath Will Accompany Any Assertion Messages in the Model
		InstancePath         : STRING           := "*";
		--
		-- 'X' generation control parameter for timing checks and path delay
		XOn                  : BOOLEAN          := TRUE;
		--
		-- Assertion messages generation control parameter for violation of timing checks
		MsgOn                : BOOLEAN          := TRUE;
		--
		-- VitalTimingCheck Switch
		TimingChecksOn       : BOOLEAN          := TRUE
	);
	PORT (
		CLK                 : IN      STD_ULOGIC := 'X';
		D                   : IN      STD_ULOGIC := 'X';
		E                   : IN      STD_ULOGIC := 'X';
		M                   : IN      STD_ULOGIC := 'X';
		IOPCL               : IN      STD_ULOGIC := 'X';
		ODE                 : IN      STD_ULOGIC := 'X';
		PAD                 : INOUT   STD_ULOGIC := 'X';
		Y                   : OUT     STD_ULOGIC := 'X'
		
	);
	--
	attribute Vital_Level0 OF FEPTML : ENTITY IS TRUE;
	--
end FEPTML;

ARCHITECTURE VITAL_ACT OF FEPTML IS
	--
	ATTRIBUTE Vital_Level1 OF VITAL_ACT : ARCHITECTURE IS TRUE;
	--
	--
	--Internal Delay Signals - delayed be the interconnect path delay
	SIGNAL    CLK_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    D_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    E_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    M_ipd                     : STD_ULOGIC := 'U';
	SIGNAL    IOPCL_ipd                 : STD_ULOGIC := 'U';
	SIGNAL    ODE_ipd                   : STD_ULOGIC := 'U';
	SIGNAL    PAD_ipd                   : STD_ULOGIC := 'U';
	
	BEGIN
	-----------------------------------------------
	-- Input Path Delay Section
	-----------------------------------------------
	WireDelay : BLOCK
	BEGIN
		VitalWireDelay (
				OutSig             => CLK_ipd,
				InSig              => CLK,
				twire              => tipd_CLK
		);
		VitalWireDelay (
				OutSig             => D_ipd,
				InSig              => D,
				twire              => tipd_D
		);
		VitalWireDelay (
				OutSig             => E_ipd,
				InSig              => E,
				twire              => tipd_E
		);
		VitalWireDelay (
				OutSig             => M_ipd,
				InSig              => M,
				twire              => tipd_M
		);
		VitalWireDelay (
				OutSig             => IOPCL_ipd,
				InSig              => IOPCL,
				twire              => tipd_IOPCL
		);
		VitalWireDelay (
				OutSig             => ODE_ipd,
				InSig              => ODE,
				twire              => tipd_ODE
		);
		VitalWireDelay (
				OutSig             => PAD_ipd,
				InSig              => PAD,
				twire              => tipd_PAD
		);
	
	END BLOCK WireDelay;
	
	-----------------------------------------------
	-- Behavior Section
	-----------------------------------------------
	VITALBehavior : PROCESS (CLK_ipd, D_ipd, E_ipd, M_ipd, IOPCL_ipd, ODE_ipd, PAD_ipd	
	                        )
		--
		-- Variable(s) for internal use in VitalPeriodPulseCheck
		VARIABLE  CLK_PeriodData            : VitalPeriodDataType := VitalPeriodDataInit;
		VARIABLE  IOPCL_PeriodData          : VitalPeriodDataType := VitalPeriodDataInit;
		--
		-- Variable(s) for internal use in VitalRecoveryRemovalCheck
		VARIABLE  IOPCL_CLK_TimingDataRR    : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) for internal use in VitalSetupHoldCheck
		VARIABLE  D_CLK_TimingDataSH        : VitalTimingDataType := VitalTimingDataInit;
		VARIABLE  ODE_CLK_TimingDataSH      : VitalTimingDataType := VitalTimingDataInit;
		--
		-- Variable(s) used in VitalPathDelay to Store GlitchData
		VARIABLE  Y_GlitchData              : VitalGlitchDataType;
		VARIABLE  PAD_GlitchData            : VitalGlitchDataType;
		--
		-- Variable(s) generated by VitalTimingCheck violation flags and/or user
		VARIABLE  SHVF_D_CLK                : STD_ULOGIC := '0';
		VARIABLE  SHVF_ODE_CLK              : STD_ULOGIC := '0';
		VARIABLE  PDVF_CLK                  : STD_ULOGIC := '0';
		VARIABLE  PDVF_IOPCL                : STD_ULOGIC := '0';
		VARIABLE  RRVF_IOPCL_CLK            : STD_ULOGIC := '0';
		VARIABLE  Violation                 : STD_ULOGIC := 'X';
		VARIABLE  FEPTML_TABStateReg        : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		VARIABLE  LSB                       : STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to store functional result
		VARIABLE  FEPTML_TAB_Result         : STD_LOGIC_VECTOR(2 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalTruthTable to store functional result
		VARIABLE  FEPTML_TTAB_Result        : STD_LOGIC_VECTOR(1 DOWNTO 1) := (OTHERS => 'X');
		--
		-- Variable(s) used in VitalStateTable to keep track of the previous values
		--VARIABLE  PrevData_FEPTML_TAB       : STD_LOGIC_VECTOR(0 TO 5);
		VARIABLE  PrevData_FEPTML_TAB       : STD_LOGIC_VECTOR(0 TO 4);
		--
		-- Variable(s) used in VitalStateTable and VitalPropagatePathDelay
		VARIABLE  Y_zd                      : STD_ULOGIC;
		VARIABLE  PAD_zd                    : STD_ULOGIC;
		VARIABLE  D_delayed                 : STD_ULOGIC;
		VARIABLE  ODE_delayed               : STD_ULOGIC;
		--
		-- State Table : FEPTML_TAB Declaration
		CONSTANT  FEPTML_TAB : VitalStateTableType (1 to 14, 1 to 8) := (
                ( '0', '0', '-', '-', '-',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '0',  '-',  '0',  '0' ),
                ( '0', '1', '/', '1', '0',  '-',  '1',  '1' ),
                ( '0', '1', '/', '0', '-',  '0',  '0',  '0' ),
                ( '0', '1', '-', '0', '-',  '0',  '0',  '0' ),
                ( '0', '-', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '-', '-', '-', '1',  '1',  '1',  '1' ),
                ( '0', '1', '/', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '-', '1', '-',  '1',  '1',  '1' ),
                ( '0', '1', '/', '-', '1',  '-',  'S',  'S' ),
                ( '0', '1', 'F', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', 'S', '-', '-',  '-',  'S',  'S' ),
                ( '0', '1', '-', '-', '1',  '-',  'S',  'S' ),
                ( 'X', '-', '-', '-', '-',  '-',  'X',  'X' ) );
	
	BEGIN
		-----------------------------------------------
		-- Timing Check Section
		-----------------------------------------------
		IF (TimingChecksOn) THEN
			-- Perform Setup/Hold Check
			--	TestSignal : D
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_D_CLK,
				TimingData         => D_CLK_TimingDataSH,
				TestSignal         => D_ipd,
				TestSignalName     => "D",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_D_CLK_noedge_posedge,
				SetupLow           => tsetup_D_CLK_noedge_posedge,
				HoldHigh           => thold_D_CLK_noedge_posedge,
				HoldLow            => thold_D_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) OR ODE_ipd ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Setup/Hold Check
			--	TestSignal : ODE
			--	RefSignal  : CLK
			VitalSetupHoldCheck (
				Violation          => SHVF_ODE_CLK,
				TimingData         => ODE_CLK_TimingDataSH,
				TestSignal         => ODE_ipd,
				TestSignalName     => "ODE",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				SetupHigh          => tsetup_ODE_CLK_noedge_posedge,
				SetupLow           => tsetup_ODE_CLK_noedge_posedge,
				HoldHigh           => thold_ODE_CLK_noedge_posedge,
				HoldLow            => thold_ODE_CLK_noedge_posedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalSetupHoldCheck
			-- Perform Recovery/Removal Check
			--	TestSignal : IOPCL
			--	RefSignal  : CLK
			VitalRecoveryRemovalCheck (
				Violation          => RRVF_IOPCL_CLK,
				TimingData         => IOPCL_CLK_TimingDataRR,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				RefSignal          => CLK_ipd,
				RefSignalName      => "CLK",
				RefDelay           => 0 ns,
				Recovery           => trecovery_IOPCL_CLK_posedge_posedge,
				Removal            => thold_IOPCL_CLK_noedge_posedge,
				ActiveLow          => TRUE,
				CheckEnabled       => TRUE,
				RefTransition      => '/',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalRecoveryRemovalCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : CLK
			VitalPeriodPulseCheck (
				Violation          => PDVF_CLK,
				PeriodData         => CLK_PeriodData,
				TestSignal         => CLK_ipd,
				TestSignalName     => "CLK",
				TestDelay          => 0 ns,
				Period             => tperiod_CLK_posedge,
				PulseWidthHigh     => tpw_CLK_posedge,
				PulseWidthLow      => tpw_CLK_negedge,
				CheckEnabled       => TO_X01 ( ( NOT IOPCL_ipd ) ) /= '1',
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
			-- Perform Minimum and Maximum Periodicity and Pulse Check
			--TestSignal : IOPCL
			VitalPeriodPulseCheck (
				Violation          => PDVF_IOPCL,
				PeriodData         => IOPCL_PeriodData,
				TestSignal         => IOPCL_ipd,
				TestSignalName     => "IOPCL",
				TestDelay          => 0 ns,
				Period             => tperiod_IOPCL,
				PulseWidthHigh     => tpw_IOPCL_posedge,
				PulseWidthLow      => tpw_IOPCL_negedge,
				CheckEnabled       => TRUE,
				HeaderMsg          => InstancePath,
				XOn                => XOn,
				MsgOn              => MsgOn,
				MsgSeverity        => WARNING
			);	--End VitalPeriodPulseCheck
		
		END IF;	--Timing Check Section
		
		-----------------------------------------------
		-- Functionality Section
		-----------------------------------------------
		

		Violation                 := PDVF_CLK or PDVF_IOPCL or RRVF_IOPCL_CLK or 
				SHVF_D_CLK or SHVF_ODE_CLK ;
		--
		--Implement Functionality for State Table : FEPTML_TAB
		VitalStateTable (
				StateTable         => FEPTML_TAB,
				--DataIn             => (Violation & IOPCL_ipd & CLK_ipd & D_ipd & ODE_ipd),
				--DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_ipd, ODE_ipd),
				DataIn             => (Violation, IOPCL_ipd, CLK_ipd, D_delayed, ODE_delayed),
				NumStates          => 1,
				Result             => FEPTML_TAB_Result,
				PreviousDataIn     => PrevData_FEPTML_TAB
		);	--End VitalStateTable
		FEPTML_TABStateReg(0)     := FEPTML_TAB_Result(2);
		LSB(0)                    := FEPTML_TAB_Result(1);
		Y_zd                      := VitalMux2(data1 => PAD_ipd, data0 => LSB(0), dselect => M_ipd);
		--
		PAD_zd := VitalBUFIF0 (data => LSB(0), enable => (NOT E_ipd));
		D_delayed := D_ipd;
		ODE_delayed := ODE_ipd;

		
		
		-----------------------------------------------
		-- Path Delay Section
		-----------------------------------------------
		VitalPathDelay01 (
				OutSignal          => Y,
				OutSignalName      => "Y",
				OutTemp            => Y_zd,
				DefaultDelay       => VitalZeroDelay01,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => PAD_ipd'LAST_EVENT,
							PathDelay       => tpd_PAD_Y,
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => tpd_IOPCL_Y,
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => M_ipd'LAST_EVENT,
							PathDelay       => tpd_M_Y,
							PathCondition   => TRUE
				                      ),
				                 3 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => tpd_CLK_Y,
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => Y_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn
		);	--End VitalPathDelay
		VitalPathDelay01Z (
				OutSignal          => PAD,
				OutSignalName      => "PAD",
				OutTemp            => PAD_zd,
				DefaultDelay       => VitalZeroDelay01Z,
				MsgSeverity        => WARNING,
				Paths              => (
				                 0 => (
							InputChangeTime => IOPCL_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_IOPCL_PAD),
							PathCondition   => TRUE
				                      ),
				                 1 => (
							InputChangeTime => CLK_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_CLK_PAD),
							PathCondition   => TRUE
				                      ),
				                 2 => (
							InputChangeTime => E_ipd'LAST_EVENT,
							PathDelay       => VitalExtendToFillDelay(tpd_E_PAD),
							PathCondition   => TRUE
				                      )
				                      ),
				GlitchData         => PAD_GlitchData,
				Mode               => OnDetect,
				XOn                => XOn,
				MsgOn              => MsgOn,
				OutputMap          => "UX01ZWLH-"
		);	--End VitalPathDelay
		
	END PROCESS VITALBehavior;

END VITAL_ACT;

configuration CFG_FEPTML_VITAL of FEPTML is
   for VITAL_ACT
   end for;
end CFG_FEPTML_VITAL;
----- CELL GAND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GAND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GAND2 : entity is TRUE;
end GAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of GAND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (G_ipd) AND (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GAND2_VITAL of GAND2 is
   for VITAL_ACT
   end for;
end CFG_GAND2_VITAL;


----- CELL GMX4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GMX4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GMX4 : entity is TRUE;
end GMX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of GMX4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (D3_ipd, D1_ipd, D2_ipd, D0_ipd),
                  dselect => (S0_ipd, G_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_Y, TRUE),
                 2 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 3 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 4 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 5 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GMX4_VITAL of GMX4 is
   for VITAL_ACT
   end for;
end CFG_GMX4_VITAL;


----- CELL GNAND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GNAND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GNAND2 : entity is TRUE;
end GNAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of GNAND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((G_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GNAND2_VITAL of GNAND2 is
   for VITAL_ACT
   end for;
end CFG_GNAND2_VITAL;


----- CELL GND -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GND is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '0');
attribute VITAL_LEVEL0 of GND : entity is TRUE;
end GND;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of GND is
   attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Y <= '0';



end VITAL_ACT;

configuration CFG_GND_VITAL of GND is
   for VITAL_ACT
   end for;
end CFG_GND_VITAL;



----- CELL GNOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GNOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GNOR2 : entity is TRUE;
end GNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of GNOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((G_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GNOR2_VITAL of GNOR2 is
   for VITAL_ACT
   end for;
end CFG_GNOR2_VITAL;


----- CELL GOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GOR2 : entity is TRUE;
end GOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of GOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (G_ipd) OR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GOR2_VITAL of GOR2 is
   for VITAL_ACT
   end for;
end CFG_GOR2_VITAL;


----- CELL GXOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GXOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GXOR2 : entity is TRUE;
end GXOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of GXOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (G_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GXOR2_VITAL of GXOR2 is
   for VITAL_ACT
   end for;
end CFG_GXOR2_VITAL;


----- CELL HA1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1 : entity is TRUE;
end HA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of HA1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (B_ipd) AND (A_ipd);
      S_zd := (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1_VITAL of HA1 is
   for VITAL_ACT
   end for;
end CFG_HA1_VITAL;


----- CELL HA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1A : entity is TRUE;
end HA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of HA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (B_ipd) AND ((NOT A_ipd));
      S_zd := (NOT ((B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1A_VITAL of HA1A is
   for VITAL_ACT
   end for;
end CFG_HA1A_VITAL;


----- CELL HA1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1B : entity is TRUE;
end HA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of HA1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (NOT ((B_ipd) AND (A_ipd)));
      S_zd := (NOT ((B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1B_VITAL of HA1B is
   for VITAL_ACT
   end for;
end CFG_HA1B_VITAL;


----- CELL HA1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1C : entity is TRUE;
end HA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of HA1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (NOT ((B_ipd) AND (A_ipd)));
      S_zd := (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1C_VITAL of HA1C is
   for VITAL_ACT
   end for;
end CFG_HA1C_VITAL;


----- CELL HCLKBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HCLKBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HCLKBUF : entity is TRUE;
end HCLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of HCLKBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HCLKBUF_VITAL of HCLKBUF is
   for VITAL_ACT
   end for;
end CFG_HCLKBUF_VITAL;


----- CELL IBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IBUF : entity is TRUE;
end IBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of IBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IBUF_VITAL of IBUF is
   for VITAL_ACT
   end for;
end CFG_IBUF_VITAL;


----- CELL INBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INBUF : entity is TRUE;
end INBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of INBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INBUF_VITAL of INBUF is
   for VITAL_ACT
   end for;
end CFG_INBUF_VITAL;


----- CELL INV -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV : entity is TRUE;
end INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of INV is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INV_VITAL of INV is
   for VITAL_ACT
   end for;
end CFG_INV_VITAL;


----- CELL INVA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INVA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INVA : entity is TRUE;
end INVA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of INVA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INVA_VITAL of INVA is
   for VITAL_ACT
   end for;
end CFG_INVA_VITAL;


----- CELL IOCLKBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IOCLKBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOCLKBUF : entity is TRUE;
end IOCLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of IOCLKBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IOCLKBUF_VITAL of IOCLKBUF is
   for VITAL_ACT
   end for;
end CFG_IOCLKBUF_VITAL;


----- CELL IODFE -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IODFE is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IODFE : entity is TRUE;
end IODFE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of IODFE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK,
          SetupLow                => tsetup_D_CLK,
          HoldHigh                => thold_D_CLK,
          HoldLow                 => thold_D_CLK,
          CheckEnabled            => 
                           TO_X01 ( E_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK,
          SetupLow                => tsetup_E_CLK,
          HoldHigh                => thold_E_CLK,
          HoldLow                 => thold_E_CLK,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IODFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IODFE_VITAL of IODFE is
   for VITAL_ACT
   end for;
end CFG_IODFE_VITAL;


----- CELL IODFEC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IODFEC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IODFEC : entity is TRUE;
end IODFEC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of IODFEC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, IOPCL_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR E_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/IODFEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_IOPCL_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IODFEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Tviol_IOPCL_CLK_posedge or Pviol_IOPCL or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               IOPCL_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (IOPCL_ipd'last_event, tpd_IOPCL_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IODFEC_VITAL of IODFEC is
   for VITAL_ACT
   end for;
end CFG_IODFEC_VITAL;


----- CELL IODFEP -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IODFEP is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IODFEP : entity is TRUE;
end IODFEP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of IODFEP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, IOPCL_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT IODFEP_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  x,  H ),
    ( x,  x,  x,  x,  H,  L,  x,  S ),
    ( x,  H,  x,  x,  U,  x,  x,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR E_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFEP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFEP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IODFEP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/IODFEP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_IOPCL_negedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IODFEP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Tviol_IOPCL_CLK_posedge or Pviol_IOPCL or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => IODFEP_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, IOPCL_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (IOPCL_ipd'last_event, tpd_IOPCL_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IODFEP_VITAL of IODFEP is
   for VITAL_ACT
   end for;
end CFG_IODFEP_VITAL;


----- CELL IOPCLBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IOPCLBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPCLBUF : entity is TRUE;
end IOPCLBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of IOPCLBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IOPCLBUF_VITAL of IOPCLBUF is
   for VITAL_ACT
   end for;
end CFG_IOPCLBUF_VITAL;


----- CELL IREC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IREC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_IDE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_IDE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      PAD                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IREC : entity is TRUE;
end IREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of IREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IDE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (IDE_ipd, IDE, tipd_IDE);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_ipd, IDE_ipd, IOPCL_ipd, PAD_ipd)

   -- timing check results
   VARIABLE Tviol_IDE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IDE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PAD_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PAD_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE IDE_delayed : STD_ULOGIC := 'X';
   VARIABLE PAD_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_IDE_CLK_posedge,
          TimingData              => Tmkr_IDE_CLK_posedge,
          TestSignal              => IDE_ipd,
          TestSignalName          => "IDE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_IDE_CLK_noedge_posedge,
          SetupLow                => tsetup_IDE_CLK_noedge_posedge,
          HoldHigh                => thold_IDE_CLK_noedge_posedge,
          HoldLow                 => thold_IDE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IREC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IREC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_PAD_CLK_posedge,
          TimingData              => Tmkr_PAD_CLK_posedge,
          TestSignal              => PAD_ipd,
          TestSignalName          => "PAD",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_PAD_CLK_noedge_posedge,
          SetupLow                => tsetup_PAD_CLK_noedge_posedge,
          HoldHigh                => thold_PAD_CLK_noedge_posedge,
          HoldLow                 => thold_PAD_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR IDE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IREC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/IREC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_IOPCL_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IREC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_IDE_CLK_posedge or Tviol_IOPCL_CLK_posedge or Tviol_PAD_CLK_posedge or Pviol_IOPCL or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               IOPCL_ipd, CLK_delayed, Q_zd, PAD_delayed, IDE_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      CLK_delayed := CLK_ipd;
      IDE_delayed := IDE_ipd;
      PAD_delayed := PAD_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (IOPCL_ipd'last_event, tpd_IOPCL_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IREC_VITAL of IREC is
   for VITAL_ACT
   end for;
end CFG_IREC_VITAL;


----- CELL IREP -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IREP is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_Q                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_IDE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_IDE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IDE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      IDE                            :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      PAD                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IREP : entity is TRUE;
end IREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of IREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IDE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (IDE_ipd, IDE, tipd_IDE);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_ipd, IDE_ipd, IOPCL_ipd, PAD_ipd)

   -- timing check results
   VARIABLE Tviol_IDE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IDE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PAD_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PAD_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE IDE_delayed : STD_ULOGIC := 'X';
   VARIABLE PAD_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_IDE_CLK_posedge,
          TimingData              => Tmkr_IDE_CLK_posedge,
          TestSignal              => IDE_ipd,
          TestSignalName          => "IDE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_IDE_CLK_noedge_posedge,
          SetupLow                => tsetup_IDE_CLK_noedge_posedge,
          HoldHigh                => thold_IDE_CLK_noedge_posedge,
          HoldLow                 => thold_IDE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IREP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IREP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_PAD_CLK_posedge,
          TimingData              => Tmkr_PAD_CLK_posedge,
          TestSignal              => PAD_ipd,
          TestSignalName          => "PAD",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_PAD_CLK_noedge_posedge,
          SetupLow                => tsetup_PAD_CLK_noedge_posedge,
          HoldHigh                => thold_PAD_CLK_noedge_posedge,
          HoldLow                 => thold_PAD_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR IDE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IREP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/IREP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_IOPCL_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IREP",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_IDE_CLK_posedge or Tviol_IOPCL_CLK_posedge or Tviol_PAD_CLK_posedge or Pviol_IOPCL or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => IODFEP_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, PAD_delayed, IDE_delayed, IOPCL_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      CLK_delayed := CLK_ipd;
      IDE_delayed := IDE_ipd;
      PAD_delayed := PAD_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (IOPCL_ipd'last_event, tpd_IOPCL_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IREP_VITAL of IREP is
   for VITAL_ACT
   end for;
end CFG_IREP_VITAL;


----- CELL JKF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF : entity is TRUE;
end JKF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of JKF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_posedge,
          TimingData              => Tmkr_J_CLK_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_posedge,
          TimingData              => Tmkr_K_CLK_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_posedge or Tviol_K_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF_VITAL of JKF is
   for VITAL_ACT
   end for;
end CFG_JKF_VITAL;


----- CELL JKF1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF1B : entity is TRUE;
end JKF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of JKF1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_negedge,
          TimingData              => Tmkr_J_CLK_negedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_negedge,
          SetupLow                => tsetup_J_CLK_noedge_negedge,
          HoldHigh                => thold_J_CLK_noedge_negedge,
          HoldLow                 => thold_J_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_negedge,
          TimingData              => Tmkr_K_CLK_negedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_negedge,
          SetupLow                => tsetup_K_CLK_noedge_negedge,
          HoldHigh                => thold_K_CLK_noedge_negedge,
          HoldLow                 => thold_K_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_negedge or Tviol_K_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF1B_VITAL of JKF1B is
   for VITAL_ACT
   end for;
end CFG_JKF1B_VITAL;


----- CELL JKF2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2A : entity is TRUE;
end JKF2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_posedge,
          TimingData              => Tmkr_J_CLK_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_posedge,
          TimingData              => Tmkr_K_CLK_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_K_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2A_VITAL of JKF2A is
   for VITAL_ACT
   end for;
end CFG_JKF2A_VITAL;


----- CELL JKF2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2B : entity is TRUE;
end JKF2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_negedge,
          TimingData              => Tmkr_J_CLK_negedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_negedge,
          SetupLow                => tsetup_J_CLK_noedge_negedge,
          HoldHigh                => thold_J_CLK_noedge_negedge,
          HoldLow                 => thold_J_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_negedge,
          TimingData              => Tmkr_K_CLK_negedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_negedge,
          SetupLow                => tsetup_K_CLK_noedge_negedge,
          HoldHigh                => thold_K_CLK_noedge_negedge,
          HoldLow                 => thold_K_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_negedge or Tviol_K_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2B_VITAL of JKF2B is
   for VITAL_ACT
   end for;
end CFG_JKF2B_VITAL;


----- CELL JKF2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2C : entity is TRUE;
end JKF2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  U,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_posedge,
          TimingData              => Tmkr_J_CLK_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_posedge,
          TimingData              => Tmkr_K_CLK_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_K_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2C_VITAL of JKF2C is
   for VITAL_ACT
   end for;
end CFG_JKF2C_VITAL;


----- CELL JKF2D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2D : entity is TRUE;
end JKF2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  U,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_negedge,
          TimingData              => Tmkr_J_CLK_negedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_negedge,
          SetupLow                => tsetup_J_CLK_noedge_negedge,
          HoldHigh                => thold_J_CLK_noedge_negedge,
          HoldLow                 => thold_J_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_negedge,
          TimingData              => Tmkr_K_CLK_negedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_negedge,
          SetupLow                => tsetup_K_CLK_noedge_negedge,
          HoldHigh                => thold_K_CLK_noedge_negedge,
          HoldLow                 => thold_K_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_negedge or Tviol_K_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2D_VITAL of JKF2D is
   for VITAL_ACT
   end for;
end CFG_JKF2D_VITAL;


----- CELL MAJ3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MAJ3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MAJ3 : entity is TRUE;
end MAJ3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of MAJ3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((C_ipd) AND (B_ipd)) OR ((B_ipd) AND (A_ipd)) OR ((C_ipd) AND
         (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MAJ3_VITAL of MAJ3 is
   for VITAL_ACT
   end for;
end CFG_MAJ3_VITAL;


----- CELL MX2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2 : entity is TRUE;
end MX2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of MX2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2_VITAL of MX2 is
   for VITAL_ACT
   end for;
end CFG_MX2_VITAL;


----- CELL MX2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2A : entity is TRUE;
end MX2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MX2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((S_ipd) AND (B_ipd)) OR (((NOT S_ipd)) AND ((NOT A_ipd))) OR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2A_VITAL of MX2A is
   for VITAL_ACT
   end for;
end CFG_MX2A_VITAL;


----- CELL MX2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2B : entity is TRUE;
end MX2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MX2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((S_ipd) AND ((NOT B_ipd))) OR (((NOT S_ipd)) AND (A_ipd)) OR ((A_ipd) AND ((NOT B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2B_VITAL of MX2B is
   for VITAL_ACT
   end for;
end CFG_MX2B_VITAL;


----- CELL MX2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2C : entity is TRUE;
end MX2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of MX2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));
      Y_zd := NOT Y_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2C_VITAL of MX2C is
   for VITAL_ACT
   end for;
end CFG_MX2C_VITAL;


----- CELL MX4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX4 : entity is TRUE;
end MX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of MX4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (D3_ipd, D2_ipd, D1_ipd, D0_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S1_ipd'last_event, tpd_S1_Y, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_Y, TRUE),
                 2 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 3 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 4 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 5 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX4_VITAL of MX4 is
   for VITAL_ACT
   end for;
end CFG_MX4_VITAL;


----- CELL MXC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MXC1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MXC1 : entity is TRUE;
end MXC1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MXC1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE MUX_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((D_ipd) AND (((B_ipd) AND (S_ipd)) OR ((A_ipd) AND ((NOT S_ipd)))))
      --   OR ((C_ipd) AND ((NOT (((B_ipd) AND (S_ipd)) OR ((A_ipd) AND ((NOT
      --   S_ipd)))))));
      MUX_Out := VitalMUX2(B_ipd, A_ipd, S_ipd);
      Y_zd := VitalMUX2(D_ipd, C_ipd, MUX_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MXC1_VITAL of MXC1 is
   for VITAL_ACT
   end for;
end CFG_MXC1_VITAL;


----- CELL MXT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MXT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0B_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0A_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0A                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0B                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0A                            :	in    STD_ULOGIC;
      S0B                            :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MXT : entity is TRUE;
end MXT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MXT is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0A_ipd, S0A, tipd_S0A);
   VitalWireDelay (S0B_ipd, S0B, tipd_S0B);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0A_ipd, S0B_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE MUX1_Out, MUX2_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((S0A_ipd) AND ((NOT S1_ipd)) AND (D1_ipd)) OR (((NOT S0A_ipd)) AND
      --   ((NOT S1_ipd)) AND (D0_ipd)) OR (((NOT S0B_ipd)) AND (S1_ipd) AND
      --   (D2_ipd)) OR ((S0B_ipd) AND (S1_ipd) AND (D3_ipd));
      MUX1_Out := VitalMUX2(D1_ipd, D0_ipd, S0A_ipd);
      MUX2_Out := VitalMUX2(D3_ipd, D2_ipd, S0B_ipd);
      Y_zd := VitalMUX2(MUX2_Out, MUX1_Out, S1_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S1_ipd'last_event, tpd_S1_Y, TRUE),
                 1 => (S0B_ipd'last_event, tpd_S0B_Y, TRUE),
                 2 => (S0A_ipd'last_event, tpd_S0A_Y, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 4 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 5 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 6 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MXT_VITAL of MXT is
   for VITAL_ACT
   end for;
end CFG_MXT_VITAL;


----- CELL NAND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND2 : entity is TRUE;
end NAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND2_VITAL of NAND2 is
   for VITAL_ACT
   end for;
end CFG_NAND2_VITAL;


----- CELL NAND2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND2A : entity is TRUE;
end NAND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND2A_VITAL of NAND2A is
   for VITAL_ACT
   end for;
end CFG_NAND2A_VITAL;


----- CELL NAND2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND2B : entity is TRUE;
end NAND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) AND ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND2B_VITAL of NAND2B is
   for VITAL_ACT
   end for;
end CFG_NAND2B_VITAL;


----- CELL NAND3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3 : entity is TRUE;
end NAND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND (A_ipd) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3_VITAL of NAND3 is
   for VITAL_ACT
   end for;
end CFG_NAND3_VITAL;


----- CELL NAND3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3A : entity is TRUE;
end NAND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND ((NOT A_ipd)) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3A_VITAL of NAND3A is
   for VITAL_ACT
   end for;
end CFG_NAND3A_VITAL;


----- CELL NAND3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3B : entity is TRUE;
end NAND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3B_VITAL of NAND3B is
   for VITAL_ACT
   end for;
end CFG_NAND3B_VITAL;


----- CELL NAND3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3C : entity is TRUE;
end NAND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3C_VITAL of NAND3C is
   for VITAL_ACT
   end for;
end CFG_NAND3C_VITAL;


----- CELL NAND4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4 : entity is TRUE;
end NAND4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND (A_ipd) AND (C_ipd) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4_VITAL of NAND4 is
   for VITAL_ACT
   end for;
end CFG_NAND4_VITAL;


----- CELL NAND4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4A : entity is TRUE;
end NAND4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4A_VITAL of NAND4A is
   for VITAL_ACT
   end for;
end CFG_NAND4A_VITAL;


----- CELL NAND4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4B : entity is TRUE;
end NAND4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4B_VITAL of NAND4B is
   for VITAL_ACT
   end for;
end CFG_NAND4B_VITAL;


----- CELL NAND4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4C : entity is TRUE;
end NAND4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4C_VITAL of NAND4C is
   for VITAL_ACT
   end for;
end CFG_NAND4C_VITAL;


----- CELL NAND4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4D : entity is TRUE;
end NAND4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND ((NOT
         D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4D_VITAL of NAND4D is
   for VITAL_ACT
   end for;
end CFG_NAND4D_VITAL;


----- CELL NAND5C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND5C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND5C : entity is TRUE;
end NAND5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NAND5C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND (D_ipd)
         AND (E_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND5C_VITAL of NAND5C is
   for VITAL_ACT
   end for;
end CFG_NAND5C_VITAL;


----- CELL NOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR2 : entity is TRUE;
end NOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR2_VITAL of NOR2 is
   for VITAL_ACT
   end for;
end CFG_NOR2_VITAL;


----- CELL NOR2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR2A : entity is TRUE;
end NOR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR2A_VITAL of NOR2A is
   for VITAL_ACT
   end for;
end CFG_NOR2A_VITAL;


----- CELL NOR2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR2B : entity is TRUE;
end NOR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) OR ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR2B_VITAL of NOR2B is
   for VITAL_ACT
   end for;
end CFG_NOR2B_VITAL;


----- CELL NOR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3 : entity is TRUE;
end NOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR (A_ipd) OR (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3_VITAL of NOR3 is
   for VITAL_ACT
   end for;
end CFG_NOR3_VITAL;


----- CELL NOR3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3A : entity is TRUE;
end NOR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR ((NOT A_ipd)) OR (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3A_VITAL of NOR3A is
   for VITAL_ACT
   end for;
end CFG_NOR3A_VITAL;


----- CELL NOR3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3B : entity is TRUE;
end NOR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3B_VITAL of NOR3B is
   for VITAL_ACT
   end for;
end CFG_NOR3B_VITAL;


----- CELL NOR3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3C : entity is TRUE;
end NOR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3C_VITAL of NOR3C is
   for VITAL_ACT
   end for;
end CFG_NOR3C_VITAL;


----- CELL NOR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4 : entity is TRUE;
end NOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR (A_ipd) OR (C_ipd) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4_VITAL of NOR4 is
   for VITAL_ACT
   end for;
end CFG_NOR4_VITAL;


----- CELL NOR4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4A : entity is TRUE;
end NOR4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4A_VITAL of NOR4A is
   for VITAL_ACT
   end for;
end CFG_NOR4A_VITAL;


----- CELL NOR4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4B : entity is TRUE;
end NOR4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4B_VITAL of NOR4B is
   for VITAL_ACT
   end for;
end CFG_NOR4B_VITAL;


----- CELL NOR4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4C : entity is TRUE;
end NOR4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4C_VITAL of NOR4C is
   for VITAL_ACT
   end for;
end CFG_NOR4C_VITAL;


----- CELL NOR4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4D : entity is TRUE;
end NOR4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR ((NOT
         D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4D_VITAL of NOR4D is
   for VITAL_ACT
   end for;
end CFG_NOR4D_VITAL;


----- CELL NOR5C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR5C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR5C : entity is TRUE;
end NOR5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of NOR5C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR (D_ipd) OR
         (E_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR5C_VITAL of NOR5C is
   for VITAL_ACT
   end for;
end CFG_NOR5C_VITAL;


----- CELL OA1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1 : entity is TRUE;
end OA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) OR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1_VITAL of OA1 is
   for VITAL_ACT
   end for;
end CFG_OA1_VITAL;


----- CELL OA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1A : entity is TRUE;
end OA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) OR ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1A_VITAL of OA1A is
   for VITAL_ACT
   end for;
end CFG_OA1A_VITAL;


----- CELL OA1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1B : entity is TRUE;
end OA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1B_VITAL of OA1B is
   for VITAL_ACT
   end for;
end CFG_OA1B_VITAL;


----- CELL OA1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1C : entity is TRUE;
end OA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1C_VITAL of OA1C is
   for VITAL_ACT
   end for;
end CFG_OA1C_VITAL;


----- CELL OA2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA2 : entity is TRUE;
end OA2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (C_ipd)) AND ((B_ipd) OR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA2_VITAL of OA2 is
   for VITAL_ACT
   end for;
end CFG_OA2_VITAL;


----- CELL OA2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA2A : entity is TRUE;
end OA2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (C_ipd)) AND ((B_ipd) OR ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA2A_VITAL of OA2A is
   for VITAL_ACT
   end for;
end CFG_OA2A_VITAL;


----- CELL OA3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA3 : entity is TRUE;
end OA3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) OR (A_ipd)) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA3_VITAL of OA3 is
   for VITAL_ACT
   end for;
end CFG_OA3_VITAL;


----- CELL OA3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA3A : entity is TRUE;
end OA3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR (A_ipd)) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA3A_VITAL of OA3A is
   for VITAL_ACT
   end for;
end CFG_OA3A_VITAL;


----- CELL OA3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA3B : entity is TRUE;
end OA3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR ((NOT A_ipd))) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA3B_VITAL of OA3B is
   for VITAL_ACT
   end for;
end CFG_OA3B_VITAL;


----- CELL OA4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA4 : entity is TRUE;
end OA4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) AND ((B_ipd) OR (A_ipd) OR (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA4_VITAL of OA4 is
   for VITAL_ACT
   end for;
end CFG_OA4_VITAL;


----- CELL OA4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA4A : entity is TRUE;
end OA4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) AND ((B_ipd) OR (A_ipd) OR ((NOT C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA4A_VITAL of OA4A is
   for VITAL_ACT
   end for;
end CFG_OA4A_VITAL;


----- CELL OA5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA5 : entity is TRUE;
end OA5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OA5 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (A_ipd)) AND ((B_ipd) OR (A_ipd) OR (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA5_VITAL of OA5 is
   for VITAL_ACT
   end for;
end CFG_OA5_VITAL;


----- CELL OAI1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI1 : entity is TRUE;
end OAI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OAI1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) AND ((B_ipd) OR (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI1_VITAL of OAI1 is
   for VITAL_ACT
   end for;
end CFG_OAI1_VITAL;


----- CELL OAI2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI2A : entity is TRUE;
end OAI2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OAI2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT D_ipd)) AND ((B_ipd) OR (A_ipd) OR (C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI2A_VITAL of OAI2A is
   for VITAL_ACT
   end for;
end CFG_OAI2A_VITAL;


----- CELL OAI3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI3 : entity is TRUE;
end OAI3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OAI3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) AND ((B_ipd) OR (A_ipd)) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI3_VITAL of OAI3 is
   for VITAL_ACT
   end for;
end CFG_OAI3_VITAL;


----- CELL OAI3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI3A : entity is TRUE;
end OAI3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OAI3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT C_ipd)) AND ((B_ipd) OR (A_ipd)) AND ((NOT D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI3A_VITAL of OAI3A is
   for VITAL_ACT
   end for;
end CFG_OAI3A_VITAL;


----- CELL OBHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OBHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OBHS : entity is TRUE;
end OBHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OBHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := TO_X01(D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OBHS_VITAL of OBHS is
   for VITAL_ACT
   end for;
end CFG_OBHS_VITAL;


----- CELL OBUFTH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OBUFTH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OBUFTH : entity is TRUE;
end OBUFTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OBUFTH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_OBUFTH_VITAL of OBUFTH is
   for VITAL_ACT
   end for;
end CFG_OBUFTH_VITAL;


----- CELL OBUFTL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OBUFTL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OBUFTL : entity is TRUE;
end OBUFTL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OBUFTL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_OBUFTL_VITAL of OBUFTL is
   for VITAL_ACT
   end for;
end CFG_OBUFTL_VITAL;


----- CELL OR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR2 : entity is TRUE;
end OR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR2_VITAL of OR2 is
   for VITAL_ACT
   end for;
end CFG_OR2_VITAL;


----- CELL OR2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR2A : entity is TRUE;
end OR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR2A_VITAL of OR2A is
   for VITAL_ACT
   end for;
end CFG_OR2A_VITAL;


----- CELL OR2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR2B : entity is TRUE;
end OR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR2B_VITAL of OR2B is
   for VITAL_ACT
   end for;
end CFG_OR2B_VITAL;


----- CELL OR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3 : entity is TRUE;
end OR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR (A_ipd) OR (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3_VITAL of OR3 is
   for VITAL_ACT
   end for;
end CFG_OR3_VITAL;


----- CELL OR3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3A : entity is TRUE;
end OR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR ((NOT A_ipd)) OR (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3A_VITAL of OR3A is
   for VITAL_ACT
   end for;
end CFG_OR3A_VITAL;


----- CELL OR3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3B : entity is TRUE;
end OR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3B_VITAL of OR3B is
   for VITAL_ACT
   end for;
end CFG_OR3B_VITAL;


----- CELL OR3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3C : entity is TRUE;
end OR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3C_VITAL of OR3C is
   for VITAL_ACT
   end for;
end CFG_OR3C_VITAL;


----- CELL OR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4 : entity is TRUE;
end OR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR (A_ipd) OR (C_ipd) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4_VITAL of OR4 is
   for VITAL_ACT
   end for;
end CFG_OR4_VITAL;


----- CELL OR4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4A : entity is TRUE;
end OR4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4A_VITAL of OR4A is
   for VITAL_ACT
   end for;
end CFG_OR4A_VITAL;


----- CELL OR4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4B : entity is TRUE;
end OR4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4B_VITAL of OR4B is
   for VITAL_ACT
   end for;
end CFG_OR4B_VITAL;


----- CELL OR4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4C : entity is TRUE;
end OR4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4C_VITAL of OR4C is
   for VITAL_ACT
   end for;
end CFG_OR4C_VITAL;


----- CELL OR4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4D : entity is TRUE;
end OR4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR ((NOT D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4D_VITAL of OR4D is
   for VITAL_ACT
   end for;
end CFG_OR4D_VITAL;


----- CELL OR5B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR5B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR5B : entity is TRUE;
end OR5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OR5B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR5B_VITAL of OR5B is
   for VITAL_ACT
   end for;
end CFG_OR5B_VITAL;


----- CELL ORECTH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ORECTH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ORECTH : entity is TRUE;
end ORECTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of ORECTH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';
   SIGNAL ODE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   VitalWireDelay (ODE_ipd, ODE, tipd_ODE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_ODE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_ODE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE ODE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zdi : STD_LOGIC is Results(1);
   VARIABLE PAD_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR ODE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORECTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORECTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_ODE_CLK_posedge,
          TimingData              => Tmkr_ODE_CLK_posedge,
          TestSignal              => ODE_ipd,
          TestSignalName          => "ODE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_ODE_CLK_noedge_posedge,
          SetupLow                => tsetup_ODE_CLK_noedge_posedge,
          HoldHigh                => thold_ODE_CLK_noedge_posedge,
          HoldLow                 => thold_ODE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORECTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/ORECTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_IOPCL_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/ORECTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_IOPCL_CLK_posedge or Pviol_IOPCL or Tviol_ODE_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zdi,
        PreviousDataIn => PrevData_PAD,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               IOPCL_ipd, CLK_delayed, PAD_zdi, D_delayed, ODE_delayed, CLK_ipd));
      PAD_zdi := Violation XOR PAD_zdi;
      PAD_zd := VitalBUFIF0 (data => PAD_zdi,
             enable => (NOT E_ipd));
      CLK_delayed := CLK_ipd;
      D_delayed := D_ipd;
      ODE_delayed := ODE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (IOPCL_ipd'last_event, VitalExtendToFillDelay(tpd_IOPCL_PAD), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 2 => (CLK_ipd'last_event, VitalExtendToFillDelay(tpd_CLK_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_ORECTH_VITAL of ORECTH is
   for VITAL_ACT
   end for;
end CFG_ORECTH_VITAL;


----- CELL ORECTL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ORECTL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ORECTL : entity is TRUE;
end ORECTL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of ORECTL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';
   SIGNAL ODE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   VitalWireDelay (ODE_ipd, ODE, tipd_ODE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_ODE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_ODE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE ODE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zdi : STD_LOGIC is Results(1);
   VARIABLE PAD_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR ODE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORECTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORECTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_ODE_CLK_posedge,
          TimingData              => Tmkr_ODE_CLK_posedge,
          TestSignal              => ODE_ipd,
          TestSignalName          => "ODE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_ODE_CLK_noedge_posedge,
          SetupLow                => tsetup_ODE_CLK_noedge_posedge,
          HoldHigh                => thold_ODE_CLK_noedge_posedge,
          HoldLow                 => thold_ODE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORECTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/ORECTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_IOPCL_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/ORECTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_IOPCL_CLK_posedge or Pviol_IOPCL or Tviol_ODE_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zdi,
        PreviousDataIn => PrevData_PAD,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               IOPCL_ipd, CLK_delayed, PAD_zdi, D_delayed, ODE_delayed, CLK_ipd));
      PAD_zdi := Violation XOR PAD_zdi;
      PAD_zd := VitalBUFIF0 (data => PAD_zdi,
             enable => (NOT E_ipd));
      CLK_delayed := CLK_ipd;
      D_delayed := D_ipd;
      ODE_delayed := ODE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (IOPCL_ipd'last_event, VitalExtendToFillDelay(tpd_IOPCL_PAD), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 2 => (CLK_ipd'last_event, VitalExtendToFillDelay(tpd_CLK_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_ORECTL_VITAL of ORECTL is
   for VITAL_ACT
   end for;
end CFG_ORECTL_VITAL;


----- CELL OREPTH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OREPTH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OREPTH : entity is TRUE;
end OREPTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of OREPTH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';
   SIGNAL ODE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   VitalWireDelay (ODE_ipd, ODE, tipd_ODE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_ODE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_ODE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE ODE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zdi : STD_LOGIC is Results(1);
   VARIABLE PAD_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT IODFEP_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  x,  H ),
    ( x,  x,  x,  x,  H,  L,  x,  S ),
    ( x,  H,  x,  x,  U,  x,  x,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR ODE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/OREPTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/OREPTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_ODE_CLK_posedge,
          TimingData              => Tmkr_ODE_CLK_posedge,
          TestSignal              => ODE_ipd,
          TestSignalName          => "ODE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_ODE_CLK_noedge_posedge,
          SetupLow                => tsetup_ODE_CLK_noedge_posedge,
          HoldHigh                => thold_ODE_CLK_noedge_posedge,
          HoldLow                 => thold_ODE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/OREPTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/OREPTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_IOPCL_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/OREPTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_IOPCL_CLK_posedge or Pviol_IOPCL or Tviol_ODE_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zdi,
        PreviousDataIn => PrevData_PAD,
        StateTable => IODFEP_Q_tab,
        DataIn => (
               CLK_delayed, PAD_zdi, D_delayed, ODE_delayed, IOPCL_ipd, CLK_ipd));
      PAD_zdi := Violation XOR PAD_zdi;
      PAD_zd := VitalBUFIF0 (data => PAD_zdi,
             enable => (NOT E_ipd));
      CLK_delayed := CLK_ipd;
      D_delayed := D_ipd;
      ODE_delayed := ODE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (IOPCL_ipd'last_event, VitalExtendToFillDelay(tpd_IOPCL_PAD), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 2 => (CLK_ipd'last_event, VitalExtendToFillDelay(tpd_CLK_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_OREPTH_VITAL of OREPTH is
   for VITAL_ACT
   end for;
end CFG_OREPTH_VITAL;


----- CELL OREPTL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OREPTL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_IOPCL_PAD                  :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_IOPCL_CLK_noedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_IOPCL_CLK_posedge_posedge            :	VitalDelayType := 0.000 ns;
      thold_ODE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_ODE_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_IOPCL_negedge              :	VitalDelayType := 0.000 ns;
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_IOPCL                     :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ODE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK                            :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      IOPCL                          :	in    STD_ULOGIC;
      ODE                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OREPTL : entity is TRUE;
end OREPTL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of OREPTL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL IOPCL_ipd	 : STD_ULOGIC := 'X';
   SIGNAL ODE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (IOPCL_ipd, IOPCL, tipd_IOPCL);
   VitalWireDelay (ODE_ipd, ODE, tipd_ODE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_ipd, D_ipd, E_ipd, IOPCL_ipd, ODE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_IOPCL_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_IOPCL_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_ODE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_ODE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_IOPCL	: STD_ULOGIC := '0';
   VARIABLE PInfo_IOPCL	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE ODE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zdi : STD_LOGIC is Results(1);
   VARIABLE PAD_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT IODFEP_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  L,  x,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  x,  H ),
    ( x,  x,  x,  x,  H,  L,  x,  S ),
    ( x,  H,  x,  x,  U,  x,  x,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) OR ODE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/OREPTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_IOPCL_CLK_posedge,
          TimingData              => Tmkr_IOPCL_CLK_posedge,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_IOPCL_CLK_posedge_posedge,
          Removal                 => thold_IOPCL_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/OREPTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_ODE_CLK_posedge,
          TimingData              => Tmkr_ODE_CLK_posedge,
          TestSignal              => ODE_ipd,
          TestSignalName          => "ODE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_ODE_CLK_noedge_posedge,
          SetupLow                => tsetup_ODE_CLK_noedge_posedge,
          HoldHigh                => thold_ODE_CLK_noedge_posedge,
          HoldLow                 => thold_ODE_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/OREPTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT IOPCL_ipd)) /= '1',
          HeaderMsg               => InstancePath &"/OREPTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_IOPCL,
          PeriodData              => PInfo_IOPCL,
          TestSignal              => IOPCL_ipd,
          TestSignalName          => "IOPCL",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_IOPCL_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/OREPTL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_IOPCL_CLK_posedge or Pviol_IOPCL or Tviol_ODE_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zdi,
        PreviousDataIn => PrevData_PAD,
        StateTable => IODFEP_Q_tab,
        DataIn => (
               CLK_delayed, PAD_zdi, D_delayed, ODE_delayed, IOPCL_ipd, CLK_ipd));
      PAD_zdi := Violation XOR PAD_zdi;
      PAD_zd := VitalBUFIF0 (data => PAD_zdi,
             enable => (NOT E_ipd));
      CLK_delayed := CLK_ipd;
      D_delayed := D_ipd;
      ODE_delayed := ODE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (IOPCL_ipd'last_event, VitalExtendToFillDelay(tpd_IOPCL_PAD), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 2 => (CLK_ipd'last_event, VitalExtendToFillDelay(tpd_CLK_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_OREPTL_VITAL of OREPTL is
   for VITAL_ACT
   end for;
end CFG_OREPTL_VITAL;


----- CELL OUTBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OUTBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OUTBUF : entity is TRUE;
end OUTBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of OUTBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := TO_X01(D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OUTBUF_VITAL of OUTBUF is
   for VITAL_ACT
   end for;
end CFG_OUTBUF_VITAL;


----- CELL TBHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TBHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TBHS : entity is TRUE;
end TBHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of TBHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_TBHS_VITAL of TBHS is
   for VITAL_ACT
   end for;
end CFG_TBHS_VITAL;


----- CELL TF1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TF1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TF1A : entity is TRUE;
end TF1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of TF1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (T_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_T_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT TF1A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( x,  L,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_posedge,
          TimingData              => Tmkr_T_CLK_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TF1A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, T_delayed, Q_zd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      T_delayed := T_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_TF1A_VITAL of TF1A is
   for VITAL_ACT
   end for;
end CFG_TF1A_VITAL;


----- CELL TF1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TF1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TF1B : entity is TRUE;
end TF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of TF1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (T_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_T_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT TF1A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( x,  L,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_negedge,
          TimingData              => Tmkr_T_CLK_negedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_T_CLK_noedge_negedge,
          SetupLow                => tsetup_T_CLK_noedge_negedge,
          HoldHigh                => thold_T_CLK_noedge_negedge,
          HoldLow                 => thold_T_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TF1A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, T_delayed, Q_zd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      T_delayed := T_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_TF1B_VITAL of TF1B is
   for VITAL_ACT
   end for;
end CFG_TF1B_VITAL;


----- CELL TRIBUFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TRIBUFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns, 0.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TRIBUFF : entity is TRUE;
end TRIBUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of TRIBUFF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_PAD), TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_TRIBUFF_VITAL of TRIBUFF is
   for VITAL_ACT
   end for;
end CFG_TRIBUFF_VITAL;


----- CELL VCC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity VCC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '1');
attribute VITAL_LEVEL0 of VCC : entity is TRUE;
end VCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of VCC is
   attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Y <= '1';



end VITAL_ACT;

configuration CFG_VCC_VITAL of VCC is
   for VITAL_ACT
   end for;
end CFG_VCC_VITAL;



----- CELL XA1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XA1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XA1 : entity is TRUE;
end XA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of XA1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) XOR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XA1_VITAL of XA1 is
   for VITAL_ACT
   end for;
end CFG_XA1_VITAL;


----- CELL XA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XA1A : entity is TRUE;
end XA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of XA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((NOT ((B_ipd) XOR (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XA1A_VITAL of XA1A is
   for VITAL_ACT
   end for;
end CFG_XA1A_VITAL;


----- CELL XNOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNOR2 : entity is TRUE;
end XNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of XNOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XNOR2_VITAL of XNOR2 is
   for VITAL_ACT
   end for;
end CFG_XNOR2_VITAL;


----- CELL XO1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XO1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XO1 : entity is TRUE;
end XO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of XO1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) XOR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XO1_VITAL of XO1 is
   for VITAL_ACT
   end for;
end CFG_XO1_VITAL;


----- CELL XO1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XO1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XO1A : entity is TRUE;
end XO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of XO1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((NOT ((B_ipd) XOR (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XO1A_VITAL of XO1A is
   for VITAL_ACT
   end for;
end CFG_XO1A_VITAL;


----- CELL XOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR2 : entity is TRUE;
end XOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library act3;
use act3.VTABLES.all;
architecture VITAL_ACT of XOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XOR2_VITAL of XOR2 is
   for VITAL_ACT
   end for;
end CFG_XOR2_VITAL;


---- end of library ----
